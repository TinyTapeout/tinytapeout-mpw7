magic
tech sky130B
magscale 1 2
timestamp 1661445026
<< metal1 >>
rect 68278 700612 68284 700664
rect 68336 700652 68342 700664
rect 105446 700652 105452 700664
rect 68336 700624 105452 700652
rect 68336 700612 68342 700624
rect 105446 700612 105452 700624
rect 105504 700612 105510 700664
rect 64138 700544 64144 700596
rect 64196 700584 64202 700596
rect 170306 700584 170312 700596
rect 64196 700556 170312 700584
rect 64196 700544 64202 700556
rect 170306 700544 170312 700556
rect 170364 700544 170370 700596
rect 36630 700476 36636 700528
rect 36688 700516 36694 700528
rect 300118 700516 300124 700528
rect 36688 700488 300124 700516
rect 36688 700476 36694 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 64230 700408 64236 700460
rect 64288 700448 64294 700460
rect 364978 700448 364984 700460
rect 64288 700420 364984 700448
rect 64288 700408 64294 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 65518 700340 65524 700392
rect 65576 700380 65582 700392
rect 429838 700380 429844 700392
rect 65576 700352 429844 700380
rect 65576 700340 65582 700352
rect 429838 700340 429844 700352
rect 429896 700340 429902 700392
rect 36538 700272 36544 700324
rect 36596 700312 36602 700324
rect 559650 700312 559656 700324
rect 36596 700284 559656 700312
rect 36596 700272 36602 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 490558 699660 490564 699712
rect 490616 699700 490622 699712
rect 494790 699700 494796 699712
rect 490616 699672 494796 699700
rect 490616 699660 490622 699672
rect 494790 699660 494796 699672
rect 494848 699660 494854 699712
rect 25682 686060 25688 686112
rect 25740 686100 25746 686112
rect 71038 686100 71044 686112
rect 25740 686072 71044 686100
rect 25740 686060 25746 686072
rect 71038 686060 71044 686072
rect 71096 686060 71102 686112
rect 212350 686060 212356 686112
rect 212408 686100 212414 686112
rect 232682 686100 232688 686112
rect 212408 686072 232688 686100
rect 212408 686060 212414 686072
rect 232682 686060 232688 686072
rect 232740 686060 232746 686112
rect 296346 686060 296352 686112
rect 296404 686100 296410 686112
rect 316770 686100 316776 686112
rect 296404 686072 316776 686100
rect 296404 686060 296410 686072
rect 316770 686060 316776 686072
rect 316828 686060 316834 686112
rect 408034 686060 408040 686112
rect 408092 686100 408098 686112
rect 428642 686100 428648 686112
rect 408092 686072 428648 686100
rect 408092 686060 408098 686072
rect 428642 686060 428648 686072
rect 428700 686060 428706 686112
rect 492030 686060 492036 686112
rect 492088 686100 492094 686112
rect 512730 686100 512736 686112
rect 492088 686072 512736 686100
rect 492088 686060 492094 686072
rect 512730 686060 512736 686072
rect 512788 686060 512794 686112
rect 36906 685992 36912 686044
rect 36964 686032 36970 686044
rect 53650 686032 53656 686044
rect 36964 686004 53656 686032
rect 36964 685992 36970 686004
rect 53650 685992 53656 686004
rect 53708 685992 53714 686044
rect 64322 685992 64328 686044
rect 64380 686032 64386 686044
rect 81434 686032 81440 686044
rect 64380 686004 81440 686032
rect 64380 685992 64386 686004
rect 81434 685992 81440 686004
rect 81492 685992 81498 686044
rect 148410 685992 148416 686044
rect 148468 686032 148474 686044
rect 165706 686032 165712 686044
rect 148468 686004 165712 686032
rect 148468 685992 148474 686004
rect 165706 685992 165712 686004
rect 165764 685992 165770 686044
rect 175458 685992 175464 686044
rect 175516 686032 175522 686044
rect 193674 686032 193680 686044
rect 175516 686004 193680 686032
rect 175516 685992 175522 686004
rect 193674 685992 193680 686004
rect 193732 685992 193738 686044
rect 203518 685992 203524 686044
rect 203576 686032 203582 686044
rect 221366 686032 221372 686044
rect 203576 686004 221372 686032
rect 203576 685992 203582 686004
rect 221366 685992 221372 686004
rect 221424 685992 221430 686044
rect 260190 685992 260196 686044
rect 260248 686032 260254 686044
rect 277670 686032 277676 686044
rect 260248 686004 277676 686032
rect 260248 685992 260254 686004
rect 277670 685992 277676 686004
rect 277728 685992 277734 686044
rect 287514 685992 287520 686044
rect 287572 686032 287578 686044
rect 305362 686032 305368 686044
rect 287572 686004 305368 686032
rect 287572 685992 287578 686004
rect 305362 685992 305368 686004
rect 305420 685992 305426 686044
rect 345658 685992 345664 686044
rect 345716 686032 345722 686044
rect 361666 686032 361672 686044
rect 345716 686004 361672 686032
rect 345716 685992 345722 686004
rect 361666 685992 361672 686004
rect 361724 685992 361730 686044
rect 371510 685992 371516 686044
rect 371568 686032 371574 686044
rect 389358 686032 389364 686044
rect 371568 686004 389364 686032
rect 371568 685992 371574 686004
rect 389358 685992 389364 686004
rect 389416 685992 389422 686044
rect 399478 685992 399484 686044
rect 399536 686032 399542 686044
rect 417694 686032 417700 686044
rect 399536 686004 417700 686032
rect 399536 685992 399542 686004
rect 417694 685992 417700 686004
rect 417752 685992 417758 686044
rect 456150 685992 456156 686044
rect 456208 686032 456214 686044
rect 473354 686032 473360 686044
rect 456208 686004 473360 686032
rect 456208 685992 456214 686004
rect 473354 685992 473360 686004
rect 473412 685992 473418 686044
rect 483474 685992 483480 686044
rect 483532 686032 483538 686044
rect 501690 686032 501696 686044
rect 483532 686004 501696 686032
rect 483532 685992 483538 686004
rect 501690 685992 501696 686004
rect 501748 685992 501754 686044
rect 36814 685924 36820 685976
rect 36872 685964 36878 685976
rect 63310 685964 63316 685976
rect 36872 685936 63316 685964
rect 36872 685924 36878 685936
rect 63310 685924 63316 685936
rect 63368 685924 63374 685976
rect 66898 685924 66904 685976
rect 66956 685964 66962 685976
rect 91094 685964 91100 685976
rect 66956 685936 91100 685964
rect 66956 685924 66962 685936
rect 91094 685924 91100 685936
rect 91152 685924 91158 685976
rect 91462 685924 91468 685976
rect 91520 685964 91526 685976
rect 109678 685964 109684 685976
rect 91520 685936 109684 685964
rect 91520 685924 91526 685936
rect 109678 685924 109684 685936
rect 109736 685924 109742 685976
rect 119430 685924 119436 685976
rect 119488 685964 119494 685976
rect 137646 685964 137652 685976
rect 119488 685936 137652 685964
rect 119488 685924 119494 685936
rect 137646 685924 137652 685936
rect 137704 685924 137710 685976
rect 156322 685924 156328 685976
rect 156380 685964 156386 685976
rect 178678 685964 178684 685976
rect 156380 685936 178684 685964
rect 156380 685924 156386 685936
rect 178678 685924 178684 685936
rect 178736 685924 178742 685976
rect 232498 685924 232504 685976
rect 232556 685964 232562 685976
rect 249702 685964 249708 685976
rect 232556 685936 249708 685964
rect 232556 685924 232562 685936
rect 249702 685924 249708 685936
rect 249760 685924 249766 685976
rect 268010 685924 268016 685976
rect 268068 685964 268074 685976
rect 287698 685964 287704 685976
rect 268068 685936 287704 685964
rect 268068 685924 268074 685936
rect 287698 685924 287704 685936
rect 287756 685924 287762 685976
rect 315482 685924 315488 685976
rect 315540 685964 315546 685976
rect 333698 685964 333704 685976
rect 315540 685936 333704 685964
rect 315540 685924 315546 685936
rect 333698 685924 333704 685936
rect 333756 685924 333762 685976
rect 352006 685924 352012 685976
rect 352064 685964 352070 685976
rect 374638 685964 374644 685976
rect 352064 685936 374644 685964
rect 352064 685924 352070 685936
rect 374638 685924 374644 685936
rect 374696 685924 374702 685976
rect 428458 685924 428464 685976
rect 428516 685964 428522 685976
rect 445662 685964 445668 685976
rect 428516 685936 445668 685964
rect 428516 685924 428522 685936
rect 445662 685924 445668 685936
rect 445720 685924 445726 685976
rect 464338 685924 464344 685976
rect 464396 685964 464402 685976
rect 483658 685964 483664 685976
rect 464396 685936 483664 685964
rect 464396 685924 464402 685936
rect 483658 685924 483664 685936
rect 483716 685924 483722 685976
rect 511442 685924 511448 685976
rect 511500 685964 511506 685976
rect 529658 685964 529664 685976
rect 511500 685936 529664 685964
rect 511500 685924 511506 685936
rect 529658 685924 529664 685936
rect 529716 685924 529722 685976
rect 542998 685924 543004 685976
rect 543056 685964 543062 685976
rect 557534 685964 557540 685976
rect 543056 685936 557540 685964
rect 543056 685924 543062 685936
rect 557534 685924 557540 685936
rect 557592 685924 557598 685976
rect 94498 685856 94504 685908
rect 94556 685896 94562 685908
rect 119338 685896 119344 685908
rect 94556 685868 119344 685896
rect 94556 685856 94562 685868
rect 119338 685856 119344 685868
rect 119396 685856 119402 685908
rect 120718 685856 120724 685908
rect 120776 685896 120782 685908
rect 147306 685896 147312 685908
rect 120776 685868 147312 685896
rect 120776 685856 120782 685868
rect 147306 685856 147312 685868
rect 147364 685856 147370 685908
rect 148318 685856 148324 685908
rect 148376 685896 148382 685908
rect 175366 685896 175372 685908
rect 148376 685868 175372 685896
rect 148376 685856 148382 685868
rect 175366 685856 175372 685868
rect 175424 685856 175430 685908
rect 177298 685856 177304 685908
rect 177356 685896 177362 685908
rect 203334 685896 203340 685908
rect 177356 685868 203340 685896
rect 177356 685856 177362 685868
rect 203334 685856 203340 685868
rect 203392 685856 203398 685908
rect 204898 685856 204904 685908
rect 204956 685896 204962 685908
rect 231026 685896 231032 685908
rect 204956 685868 231032 685896
rect 204956 685856 204962 685868
rect 231026 685856 231032 685868
rect 231084 685856 231090 685908
rect 232590 685856 232596 685908
rect 232648 685896 232654 685908
rect 259362 685896 259368 685908
rect 232648 685868 259368 685896
rect 232648 685856 232654 685868
rect 259362 685856 259368 685868
rect 259420 685856 259426 685908
rect 260098 685856 260104 685908
rect 260156 685896 260162 685908
rect 287330 685896 287336 685908
rect 260156 685868 287336 685896
rect 260156 685856 260162 685868
rect 287330 685856 287336 685868
rect 287388 685856 287394 685908
rect 289078 685856 289084 685908
rect 289136 685896 289142 685908
rect 315022 685896 315028 685908
rect 289136 685868 315028 685896
rect 289136 685856 289142 685868
rect 315022 685856 315028 685868
rect 315080 685856 315086 685908
rect 316678 685856 316684 685908
rect 316736 685896 316742 685908
rect 343358 685896 343364 685908
rect 316736 685868 343364 685896
rect 316736 685856 316742 685868
rect 343358 685856 343364 685868
rect 343416 685856 343422 685908
rect 344278 685856 344284 685908
rect 344336 685896 344342 685908
rect 371326 685896 371332 685908
rect 344336 685868 371332 685896
rect 344336 685856 344342 685868
rect 371326 685856 371332 685868
rect 371384 685856 371390 685908
rect 373258 685856 373264 685908
rect 373316 685896 373322 685908
rect 399018 685896 399024 685908
rect 373316 685868 399024 685896
rect 373316 685856 373322 685868
rect 399018 685856 399024 685868
rect 399076 685856 399082 685908
rect 400858 685856 400864 685908
rect 400916 685896 400922 685908
rect 427354 685896 427360 685908
rect 400916 685868 427360 685896
rect 400916 685856 400922 685868
rect 427354 685856 427360 685868
rect 427412 685856 427418 685908
rect 428550 685856 428556 685908
rect 428608 685896 428614 685908
rect 455322 685896 455328 685908
rect 428608 685868 455328 685896
rect 428608 685856 428614 685868
rect 455322 685856 455328 685868
rect 455380 685856 455386 685908
rect 456058 685856 456064 685908
rect 456116 685896 456122 685908
rect 483014 685896 483020 685908
rect 456116 685868 483020 685896
rect 456116 685856 456122 685868
rect 483014 685856 483020 685868
rect 483072 685856 483078 685908
rect 485038 685856 485044 685908
rect 485096 685896 485102 685908
rect 511350 685896 511356 685908
rect 485096 685868 511356 685896
rect 485096 685856 485102 685868
rect 511350 685856 511356 685868
rect 511408 685856 511414 685908
rect 512638 685856 512644 685908
rect 512696 685896 512702 685908
rect 539318 685896 539324 685908
rect 512696 685868 539324 685896
rect 512696 685856 512702 685868
rect 539318 685856 539324 685868
rect 539376 685856 539382 685908
rect 540238 685856 540244 685908
rect 540296 685896 540302 685908
rect 567194 685896 567200 685908
rect 540296 685868 567200 685896
rect 540296 685856 540302 685868
rect 567194 685856 567200 685868
rect 567252 685856 567258 685908
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 182082 683204 182088 683256
rect 182140 683244 182146 683256
rect 233234 683244 233240 683256
rect 182140 683216 233240 683244
rect 182140 683204 182146 683216
rect 233234 683204 233240 683216
rect 233292 683204 233298 683256
rect 378042 683204 378048 683256
rect 378100 683244 378106 683256
rect 429194 683244 429200 683256
rect 378100 683216 429200 683244
rect 378100 683204 378106 683216
rect 429194 683204 429200 683216
rect 429252 683204 429258 683256
rect 35618 683136 35624 683188
rect 35676 683176 35682 683188
rect 36722 683176 36728 683188
rect 35676 683148 36728 683176
rect 35676 683136 35682 683148
rect 36722 683136 36728 683148
rect 36780 683136 36786 683188
rect 42702 683136 42708 683188
rect 42760 683176 42766 683188
rect 93854 683176 93860 683188
rect 42760 683148 93860 683176
rect 42760 683136 42766 683148
rect 93854 683136 93860 683148
rect 93912 683136 93918 683188
rect 97902 683136 97908 683188
rect 97960 683176 97966 683188
rect 149054 683176 149060 683188
rect 97960 683148 149060 683176
rect 97960 683136 97966 683148
rect 149054 683136 149060 683148
rect 149112 683136 149118 683188
rect 154482 683136 154488 683188
rect 154540 683176 154546 683188
rect 205634 683176 205640 683188
rect 154540 683148 205640 683176
rect 154540 683136 154546 683148
rect 205634 683136 205640 683148
rect 205692 683136 205698 683188
rect 238662 683136 238668 683188
rect 238720 683176 238726 683188
rect 289814 683176 289820 683188
rect 238720 683148 289820 683176
rect 238720 683136 238726 683148
rect 289814 683136 289820 683148
rect 289872 683136 289878 683188
rect 293862 683136 293868 683188
rect 293920 683176 293926 683188
rect 345014 683176 345020 683188
rect 293920 683148 345020 683176
rect 293920 683136 293926 683148
rect 345014 683136 345020 683148
rect 345072 683136 345078 683188
rect 350442 683136 350448 683188
rect 350500 683176 350506 683188
rect 401594 683176 401600 683188
rect 350500 683148 401600 683176
rect 350500 683136 350506 683148
rect 401594 683136 401600 683148
rect 401652 683136 401658 683188
rect 434622 683136 434628 683188
rect 434680 683176 434686 683188
rect 485774 683176 485780 683188
rect 434680 683148 485780 683176
rect 434680 683136 434686 683148
rect 485774 683136 485780 683148
rect 485832 683136 485838 683188
rect 489822 683136 489828 683188
rect 489880 683176 489886 683188
rect 542354 683176 542360 683188
rect 489880 683148 542360 683176
rect 489880 683136 489886 683148
rect 542354 683136 542360 683148
rect 542412 683136 542418 683188
rect 541618 673820 541624 673872
rect 541676 673860 541682 673872
rect 545114 673860 545120 673872
rect 541676 673832 545120 673860
rect 541676 673820 541682 673832
rect 545114 673820 545120 673832
rect 545172 673820 545178 673872
rect 567838 670692 567844 670744
rect 567896 670732 567902 670744
rect 580166 670732 580172 670744
rect 567896 670704 580172 670732
rect 567896 670692 567902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 63586 668720 63592 668772
rect 63644 668760 63650 668772
rect 64322 668760 64328 668772
rect 63644 668732 64328 668760
rect 63644 668720 63650 668732
rect 64322 668720 64328 668732
rect 64380 668720 64386 668772
rect 147674 668720 147680 668772
rect 147732 668760 147738 668772
rect 148410 668760 148416 668772
rect 147732 668732 148416 668760
rect 147732 668720 147738 668732
rect 148410 668720 148416 668732
rect 148468 668720 148474 668772
rect 259730 668720 259736 668772
rect 259788 668760 259794 668772
rect 260190 668760 260196 668772
rect 259788 668732 260196 668760
rect 259788 668720 259794 668732
rect 260190 668720 260196 668732
rect 260248 668720 260254 668772
rect 455690 668720 455696 668772
rect 455748 668760 455754 668772
rect 456150 668760 456156 668772
rect 455748 668732 456156 668760
rect 455748 668720 455754 668732
rect 456150 668720 456156 668732
rect 456208 668720 456214 668772
rect 428642 665796 428648 665848
rect 428700 665836 428706 665848
rect 435726 665836 435732 665848
rect 428700 665808 435732 665836
rect 428700 665796 428706 665808
rect 435726 665796 435732 665808
rect 435784 665796 435790 665848
rect 287698 665456 287704 665508
rect 287756 665496 287762 665508
rect 295702 665496 295708 665508
rect 287756 665468 295708 665496
rect 287756 665456 287762 665468
rect 295702 665456 295708 665468
rect 295760 665456 295766 665508
rect 316770 665456 316776 665508
rect 316828 665496 316834 665508
rect 323670 665496 323676 665508
rect 316828 665468 323676 665496
rect 316828 665456 316834 665468
rect 323670 665456 323676 665468
rect 323728 665456 323734 665508
rect 232682 665252 232688 665304
rect 232740 665292 232746 665304
rect 239766 665292 239772 665304
rect 232740 665264 239772 665292
rect 232740 665252 232746 665264
rect 239766 665252 239772 665264
rect 239824 665252 239830 665304
rect 483658 665252 483664 665304
rect 483716 665292 483722 665304
rect 491662 665292 491668 665304
rect 483716 665264 491668 665292
rect 483716 665252 483722 665264
rect 491662 665252 491668 665264
rect 491720 665252 491726 665304
rect 512730 665252 512736 665304
rect 512788 665292 512794 665304
rect 519630 665292 519636 665304
rect 512788 665264 519636 665292
rect 512788 665252 512794 665264
rect 519630 665252 519636 665264
rect 519688 665252 519694 665304
rect 13722 665116 13728 665168
rect 13780 665156 13786 665168
rect 66254 665156 66260 665168
rect 13780 665128 66260 665156
rect 13780 665116 13786 665128
rect 66254 665116 66260 665128
rect 66312 665116 66318 665168
rect 70302 665116 70308 665168
rect 70360 665156 70366 665168
rect 121454 665156 121460 665168
rect 70360 665128 121460 665156
rect 70360 665116 70366 665128
rect 121454 665116 121460 665128
rect 121512 665116 121518 665168
rect 126882 665116 126888 665168
rect 126940 665156 126946 665168
rect 178034 665156 178040 665168
rect 126940 665128 178040 665156
rect 126940 665116 126946 665128
rect 178034 665116 178040 665128
rect 178092 665116 178098 665168
rect 209682 665116 209688 665168
rect 209740 665156 209746 665168
rect 262214 665156 262220 665168
rect 209740 665128 262220 665156
rect 209740 665116 209746 665128
rect 262214 665116 262220 665128
rect 262272 665116 262278 665168
rect 266262 665116 266268 665168
rect 266320 665156 266326 665168
rect 317414 665156 317420 665168
rect 266320 665128 317420 665156
rect 266320 665116 266326 665128
rect 317414 665116 317420 665128
rect 317472 665116 317478 665168
rect 322842 665116 322848 665168
rect 322900 665156 322906 665168
rect 373994 665156 374000 665168
rect 322900 665128 374000 665156
rect 322900 665116 322906 665128
rect 373994 665116 374000 665128
rect 374052 665116 374058 665168
rect 405642 665116 405648 665168
rect 405700 665156 405706 665168
rect 458174 665156 458180 665168
rect 405700 665128 458180 665156
rect 405700 665116 405706 665128
rect 458174 665116 458180 665128
rect 458232 665116 458238 665168
rect 462222 665116 462228 665168
rect 462280 665156 462286 665168
rect 513374 665156 513380 665168
rect 462280 665128 513380 665156
rect 462280 665116 462286 665128
rect 513374 665116 513380 665128
rect 513432 665116 513438 665168
rect 518802 665116 518808 665168
rect 518860 665156 518866 665168
rect 569954 665156 569960 665168
rect 518860 665128 569960 665156
rect 518860 665116 518866 665128
rect 569954 665116 569960 665128
rect 570012 665116 570018 665168
rect 35618 665048 35624 665100
rect 35676 665088 35682 665100
rect 36906 665088 36912 665100
rect 35676 665060 36912 665088
rect 35676 665048 35682 665060
rect 36906 665048 36912 665060
rect 36964 665048 36970 665100
rect 343542 665048 343548 665100
rect 343600 665088 343606 665100
rect 345658 665088 345664 665100
rect 343600 665060 345664 665088
rect 343600 665048 343606 665060
rect 345658 665048 345664 665060
rect 345716 665048 345722 665100
rect 71866 662328 71872 662380
rect 71924 662368 71930 662380
rect 100018 662368 100024 662380
rect 71924 662340 100024 662368
rect 71924 662328 71930 662340
rect 100018 662328 100024 662340
rect 100076 662328 100082 662380
rect 127710 662368 127716 662380
rect 103486 662340 127716 662368
rect 25682 662260 25688 662312
rect 25740 662300 25746 662312
rect 36814 662300 36820 662312
rect 25740 662272 36820 662300
rect 25740 662260 25746 662272
rect 36814 662260 36820 662272
rect 36872 662260 36878 662312
rect 42886 662260 42892 662312
rect 42944 662300 42950 662312
rect 42944 662272 45554 662300
rect 42944 662260 42950 662272
rect 15194 662192 15200 662244
rect 15252 662232 15258 662244
rect 43622 662232 43628 662244
rect 15252 662204 43628 662232
rect 15252 662192 15258 662204
rect 43622 662192 43628 662204
rect 43680 662192 43686 662244
rect 45526 662232 45554 662272
rect 53742 662260 53748 662312
rect 53800 662300 53806 662312
rect 66898 662300 66904 662312
rect 53800 662272 66904 662300
rect 53800 662260 53806 662272
rect 66898 662260 66904 662272
rect 66956 662260 66962 662312
rect 81986 662260 81992 662312
rect 82044 662300 82050 662312
rect 94498 662300 94504 662312
rect 82044 662272 94504 662300
rect 82044 662260 82050 662272
rect 94498 662260 94504 662272
rect 94556 662260 94562 662312
rect 99466 662260 99472 662312
rect 99524 662300 99530 662312
rect 103486 662300 103514 662340
rect 127710 662328 127716 662340
rect 127768 662328 127774 662380
rect 165982 662328 165988 662380
rect 166040 662368 166046 662380
rect 177298 662368 177304 662380
rect 166040 662340 177304 662368
rect 166040 662328 166046 662340
rect 177298 662328 177304 662340
rect 177356 662328 177362 662380
rect 178678 662328 178684 662380
rect 178736 662368 178742 662380
rect 184014 662368 184020 662380
rect 178736 662340 184020 662368
rect 178736 662328 178742 662340
rect 184014 662328 184020 662340
rect 184072 662328 184078 662380
rect 211706 662368 211712 662380
rect 190426 662340 211712 662368
rect 99524 662272 103514 662300
rect 99524 662260 99530 662272
rect 109678 662260 109684 662312
rect 109736 662300 109742 662312
rect 120718 662300 120724 662312
rect 109736 662272 120724 662300
rect 109736 662260 109742 662272
rect 120718 662260 120724 662272
rect 120776 662260 120782 662312
rect 137922 662260 137928 662312
rect 137980 662300 137986 662312
rect 148318 662300 148324 662312
rect 137980 662272 148324 662300
rect 137980 662260 137986 662272
rect 148318 662260 148324 662272
rect 148376 662260 148382 662312
rect 183646 662260 183652 662312
rect 183704 662300 183710 662312
rect 190426 662300 190454 662340
rect 211706 662328 211712 662340
rect 211764 662328 211770 662380
rect 277670 662328 277676 662380
rect 277728 662368 277734 662380
rect 289078 662368 289084 662380
rect 277728 662340 289084 662368
rect 277728 662328 277734 662340
rect 289078 662328 289084 662340
rect 289136 662328 289142 662380
rect 306006 662328 306012 662380
rect 306064 662368 306070 662380
rect 316678 662368 316684 662380
rect 306064 662340 316684 662368
rect 306064 662328 306070 662340
rect 316678 662328 316684 662340
rect 316736 662328 316742 662380
rect 361666 662328 361672 662380
rect 361724 662368 361730 662380
rect 373258 662368 373264 662380
rect 361724 662340 373264 662368
rect 361724 662328 361730 662340
rect 373258 662328 373264 662340
rect 373316 662328 373322 662380
rect 374638 662328 374644 662380
rect 374696 662368 374702 662380
rect 379698 662368 379704 662380
rect 374696 662340 379704 662368
rect 374696 662328 374702 662340
rect 379698 662328 379704 662340
rect 379756 662328 379762 662380
rect 408034 662368 408040 662380
rect 383626 662340 408040 662368
rect 183704 662272 190454 662300
rect 183704 662260 183710 662272
rect 193674 662260 193680 662312
rect 193732 662300 193738 662312
rect 204898 662300 204904 662312
rect 193732 662272 204904 662300
rect 193732 662260 193738 662272
rect 204898 662260 204904 662272
rect 204956 662260 204962 662312
rect 222010 662260 222016 662312
rect 222068 662300 222074 662312
rect 232590 662300 232596 662312
rect 222068 662272 232596 662300
rect 222068 662260 222074 662272
rect 232590 662260 232596 662272
rect 232648 662260 232654 662312
rect 249610 662260 249616 662312
rect 249668 662300 249674 662312
rect 260098 662300 260104 662312
rect 249668 662272 260104 662300
rect 249668 662260 249674 662272
rect 260098 662260 260104 662272
rect 260156 662260 260162 662312
rect 333882 662260 333888 662312
rect 333940 662300 333946 662312
rect 344278 662300 344284 662312
rect 333940 662272 344284 662300
rect 333940 662260 333946 662272
rect 344278 662260 344284 662272
rect 344336 662260 344342 662312
rect 379606 662260 379612 662312
rect 379664 662300 379670 662312
rect 383626 662300 383654 662340
rect 408034 662328 408040 662340
rect 408092 662328 408098 662380
rect 473998 662328 474004 662380
rect 474056 662368 474062 662380
rect 485038 662368 485044 662380
rect 474056 662340 485044 662368
rect 474056 662328 474062 662340
rect 485038 662328 485044 662340
rect 485096 662328 485102 662380
rect 501690 662328 501696 662380
rect 501748 662368 501754 662380
rect 512638 662368 512644 662380
rect 501748 662340 512644 662368
rect 501748 662328 501754 662340
rect 512638 662328 512644 662340
rect 512696 662328 512702 662380
rect 518986 662328 518992 662380
rect 519044 662368 519050 662380
rect 547874 662368 547880 662380
rect 519044 662340 547880 662368
rect 519044 662328 519050 662340
rect 547874 662328 547880 662340
rect 547932 662328 547938 662380
rect 379664 662272 383654 662300
rect 379664 662260 379670 662272
rect 390002 662260 390008 662312
rect 390060 662300 390066 662312
rect 400858 662300 400864 662312
rect 390060 662272 400864 662300
rect 390060 662260 390066 662272
rect 400858 662260 400864 662272
rect 400916 662260 400922 662312
rect 417694 662260 417700 662312
rect 417752 662300 417758 662312
rect 428550 662300 428556 662312
rect 417752 662272 428556 662300
rect 417752 662260 417758 662272
rect 428550 662260 428556 662272
rect 428608 662260 428614 662312
rect 445662 662260 445668 662312
rect 445720 662300 445726 662312
rect 456058 662300 456064 662312
rect 445720 662272 456064 662300
rect 445720 662260 445726 662272
rect 456058 662260 456064 662272
rect 456116 662260 456122 662312
rect 539318 662260 539324 662312
rect 539376 662300 539382 662312
rect 542998 662300 543004 662312
rect 539376 662272 543004 662300
rect 539376 662260 539382 662272
rect 542998 662260 543004 662272
rect 543056 662260 543062 662312
rect 71958 662232 71964 662244
rect 45526 662204 71964 662232
rect 71958 662192 71964 662204
rect 72016 662192 72022 662244
rect 127066 662192 127072 662244
rect 127124 662232 127130 662244
rect 155954 662232 155960 662244
rect 127124 662204 155960 662232
rect 127124 662192 127130 662204
rect 155954 662192 155960 662204
rect 156012 662192 156018 662244
rect 238846 662192 238852 662244
rect 238904 662232 238910 662244
rect 268010 662232 268016 662244
rect 238904 662204 268016 662232
rect 238904 662192 238910 662204
rect 268010 662192 268016 662204
rect 268068 662192 268074 662244
rect 323026 662192 323032 662244
rect 323084 662232 323090 662244
rect 352006 662232 352012 662244
rect 323084 662204 352012 662232
rect 323084 662192 323090 662204
rect 352006 662192 352012 662204
rect 352064 662192 352070 662244
rect 434806 662192 434812 662244
rect 434864 662232 434870 662244
rect 463786 662232 463792 662244
rect 434864 662204 463792 662232
rect 434864 662192 434870 662204
rect 463786 662192 463792 662204
rect 463844 662192 463850 662244
rect 529658 662192 529664 662244
rect 529716 662232 529722 662244
rect 540238 662232 540244 662244
rect 529716 662204 540244 662232
rect 529716 662192 529722 662204
rect 540238 662192 540244 662204
rect 540296 662192 540302 662244
rect 16022 658928 16028 658980
rect 16080 658968 16086 658980
rect 547874 658968 547880 658980
rect 16080 658940 547880 658968
rect 16080 658928 16086 658940
rect 547874 658928 547880 658940
rect 547932 658928 547938 658980
rect 25682 658452 25688 658504
rect 25740 658492 25746 658504
rect 66898 658492 66904 658504
rect 25740 658464 66904 658492
rect 25740 658452 25746 658464
rect 66898 658452 66904 658464
rect 66956 658452 66962 658504
rect 212350 658452 212356 658504
rect 212408 658492 212414 658504
rect 232682 658492 232688 658504
rect 212408 658464 232688 658492
rect 212408 658452 212414 658464
rect 232682 658452 232688 658464
rect 232740 658452 232746 658504
rect 296346 658452 296352 658504
rect 296404 658492 296410 658504
rect 316770 658492 316776 658504
rect 296404 658464 316776 658492
rect 296404 658452 296410 658464
rect 316770 658452 316776 658464
rect 316828 658452 316834 658504
rect 408034 658452 408040 658504
rect 408092 658492 408098 658504
rect 428642 658492 428648 658504
rect 408092 658464 428648 658492
rect 408092 658452 408098 658464
rect 428642 658452 428648 658464
rect 428700 658452 428706 658504
rect 492030 658452 492036 658504
rect 492088 658492 492094 658504
rect 512730 658492 512736 658504
rect 492088 658464 512736 658492
rect 492088 658452 492094 658464
rect 512730 658452 512736 658464
rect 512788 658452 512794 658504
rect 36998 658384 37004 658436
rect 37056 658424 37062 658436
rect 53650 658424 53656 658436
rect 37056 658396 53656 658424
rect 37056 658384 37062 658396
rect 53650 658384 53656 658396
rect 53708 658384 53714 658436
rect 148318 658384 148324 658436
rect 148376 658424 148382 658436
rect 165706 658424 165712 658436
rect 148376 658396 165712 658424
rect 148376 658384 148382 658396
rect 165706 658384 165712 658396
rect 165764 658384 165770 658436
rect 175458 658384 175464 658436
rect 175516 658424 175522 658436
rect 193674 658424 193680 658436
rect 175516 658396 193680 658424
rect 175516 658384 175522 658396
rect 193674 658384 193680 658396
rect 193732 658384 193738 658436
rect 203518 658384 203524 658436
rect 203576 658424 203582 658436
rect 221366 658424 221372 658436
rect 203576 658396 221372 658424
rect 203576 658384 203582 658396
rect 221366 658384 221372 658396
rect 221424 658384 221430 658436
rect 260190 658384 260196 658436
rect 260248 658424 260254 658436
rect 277670 658424 277676 658436
rect 260248 658396 277676 658424
rect 260248 658384 260254 658396
rect 277670 658384 277676 658396
rect 277728 658384 277734 658436
rect 287514 658384 287520 658436
rect 287572 658424 287578 658436
rect 305362 658424 305368 658436
rect 287572 658396 305368 658424
rect 287572 658384 287578 658396
rect 305362 658384 305368 658396
rect 305420 658384 305426 658436
rect 345658 658384 345664 658436
rect 345716 658424 345722 658436
rect 361666 658424 361672 658436
rect 345716 658396 361672 658424
rect 345716 658384 345722 658396
rect 361666 658384 361672 658396
rect 361724 658384 361730 658436
rect 371510 658384 371516 658436
rect 371568 658424 371574 658436
rect 389358 658424 389364 658436
rect 371568 658396 389364 658424
rect 371568 658384 371574 658396
rect 389358 658384 389364 658396
rect 389416 658384 389422 658436
rect 399478 658384 399484 658436
rect 399536 658424 399542 658436
rect 417694 658424 417700 658436
rect 399536 658396 417700 658424
rect 399536 658384 399542 658396
rect 417694 658384 417700 658396
rect 417752 658384 417758 658436
rect 456058 658384 456064 658436
rect 456116 658424 456122 658436
rect 473354 658424 473360 658436
rect 456116 658396 473360 658424
rect 456116 658384 456122 658396
rect 473354 658384 473360 658396
rect 473412 658384 473418 658436
rect 483474 658384 483480 658436
rect 483532 658424 483538 658436
rect 501690 658424 501696 658436
rect 483532 658396 501696 658424
rect 483532 658384 483538 658396
rect 501690 658384 501696 658396
rect 501748 658384 501754 658436
rect 36906 658316 36912 658368
rect 36964 658356 36970 658368
rect 63310 658356 63316 658368
rect 36964 658328 63316 658356
rect 36964 658316 36970 658328
rect 63310 658316 63316 658328
rect 63368 658316 63374 658368
rect 64322 658316 64328 658368
rect 64380 658356 64386 658368
rect 81434 658356 81440 658368
rect 64380 658328 81440 658356
rect 64380 658316 64386 658328
rect 81434 658316 81440 658328
rect 81492 658316 81498 658368
rect 91462 658316 91468 658368
rect 91520 658356 91526 658368
rect 109678 658356 109684 658368
rect 91520 658328 109684 658356
rect 91520 658316 91526 658328
rect 109678 658316 109684 658328
rect 109736 658316 109742 658368
rect 119430 658316 119436 658368
rect 119488 658356 119494 658368
rect 137646 658356 137652 658368
rect 119488 658328 137652 658356
rect 119488 658316 119494 658328
rect 137646 658316 137652 658328
rect 137704 658316 137710 658368
rect 156322 658316 156328 658368
rect 156380 658356 156386 658368
rect 178678 658356 178684 658368
rect 156380 658328 178684 658356
rect 156380 658316 156386 658328
rect 178678 658316 178684 658328
rect 178736 658316 178742 658368
rect 232590 658316 232596 658368
rect 232648 658356 232654 658368
rect 249702 658356 249708 658368
rect 232648 658328 249708 658356
rect 232648 658316 232654 658328
rect 249702 658316 249708 658328
rect 249760 658316 249766 658368
rect 268010 658316 268016 658368
rect 268068 658356 268074 658368
rect 287698 658356 287704 658368
rect 268068 658328 287704 658356
rect 268068 658316 268074 658328
rect 287698 658316 287704 658328
rect 287756 658316 287762 658368
rect 315482 658316 315488 658368
rect 315540 658356 315546 658368
rect 333698 658356 333704 658368
rect 315540 658328 333704 658356
rect 315540 658316 315546 658328
rect 333698 658316 333704 658328
rect 333756 658316 333762 658368
rect 352006 658316 352012 658368
rect 352064 658356 352070 658368
rect 374638 658356 374644 658368
rect 352064 658328 374644 658356
rect 352064 658316 352070 658328
rect 374638 658316 374644 658328
rect 374696 658316 374702 658368
rect 428458 658316 428464 658368
rect 428516 658356 428522 658368
rect 445662 658356 445668 658368
rect 428516 658328 445668 658356
rect 428516 658316 428522 658328
rect 445662 658316 445668 658328
rect 445720 658316 445726 658368
rect 464338 658316 464344 658368
rect 464396 658356 464402 658368
rect 483658 658356 483664 658368
rect 464396 658328 483664 658356
rect 464396 658316 464402 658328
rect 483658 658316 483664 658328
rect 483716 658316 483722 658368
rect 511442 658316 511448 658368
rect 511500 658356 511506 658368
rect 529658 658356 529664 658368
rect 511500 658328 529664 658356
rect 511500 658316 511506 658328
rect 529658 658316 529664 658328
rect 529716 658316 529722 658368
rect 542998 658316 543004 658368
rect 543056 658356 543062 658368
rect 557534 658356 557540 658368
rect 543056 658328 557540 658356
rect 543056 658316 543062 658328
rect 557534 658316 557540 658328
rect 557592 658316 557598 658368
rect 69658 658248 69664 658300
rect 69716 658288 69722 658300
rect 91094 658288 91100 658300
rect 69716 658260 91100 658288
rect 69716 658248 69722 658260
rect 91094 658248 91100 658260
rect 91152 658248 91158 658300
rect 94498 658248 94504 658300
rect 94556 658288 94562 658300
rect 119338 658288 119344 658300
rect 94556 658260 119344 658288
rect 94556 658248 94562 658260
rect 119338 658248 119344 658260
rect 119396 658248 119402 658300
rect 120718 658248 120724 658300
rect 120776 658288 120782 658300
rect 147306 658288 147312 658300
rect 120776 658260 147312 658288
rect 120776 658248 120782 658260
rect 147306 658248 147312 658260
rect 147364 658248 147370 658300
rect 148410 658248 148416 658300
rect 148468 658288 148474 658300
rect 175366 658288 175372 658300
rect 148468 658260 175372 658288
rect 148468 658248 148474 658260
rect 175366 658248 175372 658260
rect 175424 658248 175430 658300
rect 177298 658248 177304 658300
rect 177356 658288 177362 658300
rect 203334 658288 203340 658300
rect 177356 658260 203340 658288
rect 177356 658248 177362 658260
rect 203334 658248 203340 658260
rect 203392 658248 203398 658300
rect 204898 658248 204904 658300
rect 204956 658288 204962 658300
rect 231026 658288 231032 658300
rect 204956 658260 231032 658288
rect 204956 658248 204962 658260
rect 231026 658248 231032 658260
rect 231084 658248 231090 658300
rect 232498 658248 232504 658300
rect 232556 658288 232562 658300
rect 259362 658288 259368 658300
rect 232556 658260 259368 658288
rect 232556 658248 232562 658260
rect 259362 658248 259368 658260
rect 259420 658248 259426 658300
rect 260098 658248 260104 658300
rect 260156 658288 260162 658300
rect 287330 658288 287336 658300
rect 260156 658260 287336 658288
rect 260156 658248 260162 658260
rect 287330 658248 287336 658260
rect 287388 658248 287394 658300
rect 289078 658248 289084 658300
rect 289136 658288 289142 658300
rect 315022 658288 315028 658300
rect 289136 658260 315028 658288
rect 289136 658248 289142 658260
rect 315022 658248 315028 658260
rect 315080 658248 315086 658300
rect 316678 658248 316684 658300
rect 316736 658288 316742 658300
rect 343358 658288 343364 658300
rect 316736 658260 343364 658288
rect 316736 658248 316742 658260
rect 343358 658248 343364 658260
rect 343416 658248 343422 658300
rect 344278 658248 344284 658300
rect 344336 658288 344342 658300
rect 371326 658288 371332 658300
rect 344336 658260 371332 658288
rect 344336 658248 344342 658260
rect 371326 658248 371332 658260
rect 371384 658248 371390 658300
rect 373258 658248 373264 658300
rect 373316 658288 373322 658300
rect 399018 658288 399024 658300
rect 373316 658260 399024 658288
rect 373316 658248 373322 658260
rect 399018 658248 399024 658260
rect 399076 658248 399082 658300
rect 400858 658248 400864 658300
rect 400916 658288 400922 658300
rect 427354 658288 427360 658300
rect 400916 658260 427360 658288
rect 400916 658248 400922 658260
rect 427354 658248 427360 658260
rect 427412 658248 427418 658300
rect 428550 658248 428556 658300
rect 428608 658288 428614 658300
rect 455322 658288 455328 658300
rect 428608 658260 455328 658288
rect 428608 658248 428614 658260
rect 455322 658248 455328 658260
rect 455380 658248 455386 658300
rect 456150 658248 456156 658300
rect 456208 658288 456214 658300
rect 483014 658288 483020 658300
rect 456208 658260 483020 658288
rect 456208 658248 456214 658260
rect 483014 658248 483020 658260
rect 483072 658248 483078 658300
rect 485038 658248 485044 658300
rect 485096 658288 485102 658300
rect 511350 658288 511356 658300
rect 485096 658260 511356 658288
rect 485096 658248 485102 658260
rect 511350 658248 511356 658260
rect 511408 658248 511414 658300
rect 512638 658248 512644 658300
rect 512696 658288 512702 658300
rect 539318 658288 539324 658300
rect 512696 658260 539324 658288
rect 512696 658248 512702 658260
rect 539318 658248 539324 658260
rect 539376 658248 539382 658300
rect 540238 658248 540244 658300
rect 540296 658288 540302 658300
rect 567194 658288 567200 658300
rect 540296 658260 567200 658288
rect 540296 658248 540302 658260
rect 567194 658248 567200 658260
rect 567252 658248 567258 658300
rect 37918 657500 37924 657552
rect 37976 657540 37982 657552
rect 545758 657540 545764 657552
rect 37976 657512 545764 657540
rect 37976 657500 37982 657512
rect 545758 657500 545764 657512
rect 545816 657500 545822 657552
rect 35618 656888 35624 656940
rect 35676 656928 35682 656940
rect 36814 656928 36820 656940
rect 35676 656900 36820 656928
rect 35676 656888 35682 656900
rect 36814 656888 36820 656900
rect 36872 656888 36878 656940
rect 183554 655664 183560 655716
rect 183612 655704 183618 655716
rect 233234 655704 233240 655716
rect 183612 655676 233240 655704
rect 183612 655664 183618 655676
rect 233234 655664 233240 655676
rect 233292 655664 233298 655716
rect 378042 655664 378048 655716
rect 378100 655704 378106 655716
rect 429194 655704 429200 655716
rect 378100 655676 429200 655704
rect 378100 655664 378106 655676
rect 429194 655664 429200 655676
rect 429252 655664 429258 655716
rect 463694 655664 463700 655716
rect 463752 655704 463758 655716
rect 513374 655704 513380 655716
rect 463752 655676 513380 655704
rect 463752 655664 463758 655676
rect 513374 655664 513380 655676
rect 513432 655664 513438 655716
rect 42702 655596 42708 655648
rect 42760 655636 42766 655648
rect 93854 655636 93860 655648
rect 42760 655608 93860 655636
rect 42760 655596 42766 655608
rect 93854 655596 93860 655608
rect 93912 655596 93918 655648
rect 97902 655596 97908 655648
rect 97960 655636 97966 655648
rect 149054 655636 149060 655648
rect 97960 655608 149060 655636
rect 97960 655596 97966 655608
rect 149054 655596 149060 655608
rect 149112 655596 149118 655648
rect 154482 655596 154488 655648
rect 154540 655636 154546 655648
rect 205634 655636 205640 655648
rect 154540 655608 205640 655636
rect 154540 655596 154546 655608
rect 205634 655596 205640 655608
rect 205692 655596 205698 655648
rect 238662 655596 238668 655648
rect 238720 655636 238726 655648
rect 289814 655636 289820 655648
rect 238720 655608 289820 655636
rect 238720 655596 238726 655608
rect 289814 655596 289820 655608
rect 289872 655596 289878 655648
rect 293862 655596 293868 655648
rect 293920 655636 293926 655648
rect 345014 655636 345020 655648
rect 293920 655608 345020 655636
rect 293920 655596 293926 655608
rect 345014 655596 345020 655608
rect 345072 655596 345078 655648
rect 350442 655596 350448 655648
rect 350500 655636 350506 655648
rect 401594 655636 401600 655648
rect 350500 655608 401600 655636
rect 350500 655596 350506 655608
rect 401594 655596 401600 655608
rect 401652 655596 401658 655648
rect 434622 655596 434628 655648
rect 434680 655636 434686 655648
rect 485774 655636 485780 655648
rect 434680 655608 485780 655636
rect 434680 655596 434686 655608
rect 485774 655596 485780 655608
rect 485832 655596 485838 655648
rect 518802 655596 518808 655648
rect 518860 655636 518866 655648
rect 569954 655636 569960 655648
rect 518860 655608 569960 655636
rect 518860 655596 518866 655608
rect 569954 655596 569960 655608
rect 570012 655596 570018 655648
rect 13722 655528 13728 655580
rect 13780 655568 13786 655580
rect 66254 655568 66260 655580
rect 13780 655540 66260 655568
rect 13780 655528 13786 655540
rect 66254 655528 66260 655540
rect 66312 655528 66318 655580
rect 70302 655528 70308 655580
rect 70360 655568 70366 655580
rect 121454 655568 121460 655580
rect 70360 655540 121460 655568
rect 70360 655528 70366 655540
rect 121454 655528 121460 655540
rect 121512 655528 121518 655580
rect 126882 655528 126888 655580
rect 126940 655568 126946 655580
rect 178034 655568 178040 655580
rect 126940 655540 178040 655568
rect 126940 655528 126946 655540
rect 178034 655528 178040 655540
rect 178092 655528 178098 655580
rect 209682 655528 209688 655580
rect 209740 655568 209746 655580
rect 262214 655568 262220 655580
rect 209740 655540 262220 655568
rect 209740 655528 209746 655540
rect 262214 655528 262220 655540
rect 262272 655528 262278 655580
rect 266262 655528 266268 655580
rect 266320 655568 266326 655580
rect 317414 655568 317420 655580
rect 266320 655540 317420 655568
rect 266320 655528 266326 655540
rect 317414 655528 317420 655540
rect 317472 655528 317478 655580
rect 322842 655528 322848 655580
rect 322900 655568 322906 655580
rect 373994 655568 374000 655580
rect 322900 655540 374000 655568
rect 322900 655528 322906 655540
rect 373994 655528 374000 655540
rect 374052 655528 374058 655580
rect 405642 655528 405648 655580
rect 405700 655568 405706 655580
rect 458174 655568 458180 655580
rect 405700 655540 458180 655568
rect 405700 655528 405706 655540
rect 458174 655528 458180 655540
rect 458232 655528 458238 655580
rect 489822 655528 489828 655580
rect 489880 655568 489886 655580
rect 542354 655568 542360 655580
rect 489880 655540 542360 655568
rect 489880 655528 489886 655540
rect 542354 655528 542360 655540
rect 542412 655528 542418 655580
rect 182082 654032 182088 654084
rect 182140 654072 182146 654084
rect 183554 654072 183560 654084
rect 182140 654044 183560 654072
rect 182140 654032 182146 654044
rect 183554 654032 183560 654044
rect 183612 654032 183618 654084
rect 462222 654032 462228 654084
rect 462280 654072 462286 654084
rect 463694 654072 463700 654084
rect 462280 654044 463700 654072
rect 462280 654032 462286 654044
rect 463694 654032 463700 654044
rect 463752 654032 463758 654084
rect 63586 640772 63592 640824
rect 63644 640812 63650 640824
rect 64322 640812 64328 640824
rect 63644 640784 64328 640812
rect 63644 640772 63650 640784
rect 64322 640772 64328 640784
rect 64380 640772 64386 640824
rect 259730 640772 259736 640824
rect 259788 640812 259794 640824
rect 260190 640812 260196 640824
rect 259788 640784 260196 640812
rect 259788 640772 259794 640784
rect 260190 640772 260196 640784
rect 260248 640772 260254 640824
rect 287698 639752 287704 639804
rect 287756 639792 287762 639804
rect 295702 639792 295708 639804
rect 287756 639764 295708 639792
rect 287756 639752 287762 639764
rect 295702 639752 295708 639764
rect 295760 639752 295766 639804
rect 428642 639548 428648 639600
rect 428700 639588 428706 639600
rect 435726 639588 435732 639600
rect 428700 639560 435732 639588
rect 428700 639548 428706 639560
rect 435726 639548 435732 639560
rect 435784 639548 435790 639600
rect 232682 639344 232688 639396
rect 232740 639384 232746 639396
rect 239766 639384 239772 639396
rect 232740 639356 239772 639384
rect 232740 639344 232746 639356
rect 239766 639344 239772 639356
rect 239824 639344 239830 639396
rect 316770 639344 316776 639396
rect 316828 639384 316834 639396
rect 323670 639384 323676 639396
rect 316828 639356 323676 639384
rect 316828 639344 316834 639356
rect 323670 639344 323676 639356
rect 323728 639344 323734 639396
rect 483658 639344 483664 639396
rect 483716 639384 483722 639396
rect 491662 639384 491668 639396
rect 483716 639356 491668 639384
rect 483716 639344 483722 639356
rect 491662 639344 491668 639356
rect 491720 639344 491726 639396
rect 512730 639072 512736 639124
rect 512788 639112 512794 639124
rect 519630 639112 519636 639124
rect 512788 639084 519636 639112
rect 512788 639072 512794 639084
rect 519630 639072 519636 639084
rect 519688 639072 519694 639124
rect 35618 637508 35624 637560
rect 35676 637548 35682 637560
rect 36998 637548 37004 637560
rect 35676 637520 37004 637548
rect 35676 637508 35682 637520
rect 36998 637508 37004 637520
rect 37056 637508 37062 637560
rect 343634 637508 343640 637560
rect 343692 637548 343698 637560
rect 345658 637548 345664 637560
rect 343692 637520 345664 637548
rect 343692 637508 343698 637520
rect 345658 637508 345664 637520
rect 345716 637508 345722 637560
rect 25682 634720 25688 634772
rect 25740 634760 25746 634772
rect 36906 634760 36912 634772
rect 25740 634732 36912 634760
rect 25740 634720 25746 634732
rect 36906 634720 36912 634732
rect 36964 634720 36970 634772
rect 178678 634720 178684 634772
rect 178736 634760 178742 634772
rect 184014 634760 184020 634772
rect 178736 634732 184020 634760
rect 178736 634720 178742 634732
rect 184014 634720 184020 634732
rect 184072 634720 184078 634772
rect 231578 634720 231584 634772
rect 231636 634760 231642 634772
rect 232590 634760 232596 634772
rect 231636 634732 232596 634760
rect 231636 634720 231642 634732
rect 232590 634720 232596 634732
rect 232648 634720 232654 634772
rect 374638 634720 374644 634772
rect 374696 634760 374702 634772
rect 379698 634760 379704 634772
rect 374696 634732 379704 634760
rect 374696 634720 374702 634732
rect 379698 634720 379704 634732
rect 379756 634720 379762 634772
rect 539318 634720 539324 634772
rect 539376 634760 539382 634772
rect 542998 634760 543004 634772
rect 539376 634732 543004 634760
rect 539376 634720 539382 634732
rect 542998 634720 543004 634732
rect 543056 634720 543062 634772
rect 15194 634652 15200 634704
rect 15252 634692 15258 634704
rect 43990 634692 43996 634704
rect 15252 634664 43996 634692
rect 15252 634652 15258 634664
rect 43990 634652 43996 634664
rect 44048 634652 44054 634704
rect 71038 634652 71044 634704
rect 71096 634692 71102 634704
rect 567194 634692 567200 634704
rect 71096 634664 567200 634692
rect 71096 634652 71102 634664
rect 567194 634652 567200 634664
rect 567252 634652 567258 634704
rect 53650 634584 53656 634636
rect 53708 634624 53714 634636
rect 69658 634624 69664 634636
rect 53708 634596 69664 634624
rect 53708 634584 53714 634596
rect 69658 634584 69664 634596
rect 69716 634584 69722 634636
rect 71866 634584 71872 634636
rect 71924 634624 71930 634636
rect 100018 634624 100024 634636
rect 71924 634596 100024 634624
rect 71924 634584 71930 634596
rect 100018 634584 100024 634596
rect 100076 634584 100082 634636
rect 127986 634624 127992 634636
rect 103486 634596 127992 634624
rect 42886 634516 42892 634568
rect 42944 634556 42950 634568
rect 71958 634556 71964 634568
rect 42944 634528 71964 634556
rect 42944 634516 42950 634528
rect 71958 634516 71964 634528
rect 72016 634516 72022 634568
rect 81986 634516 81992 634568
rect 82044 634556 82050 634568
rect 94498 634556 94504 634568
rect 82044 634528 94504 634556
rect 82044 634516 82050 634528
rect 94498 634516 94504 634528
rect 94556 634516 94562 634568
rect 99466 634516 99472 634568
rect 99524 634556 99530 634568
rect 103486 634556 103514 634596
rect 127986 634584 127992 634596
rect 128044 634584 128050 634636
rect 155954 634624 155960 634636
rect 132466 634596 155960 634624
rect 99524 634528 103514 634556
rect 99524 634516 99530 634528
rect 109678 634516 109684 634568
rect 109736 634556 109742 634568
rect 120718 634556 120724 634568
rect 109736 634528 120724 634556
rect 109736 634516 109742 634528
rect 120718 634516 120724 634528
rect 120776 634516 120782 634568
rect 127066 634516 127072 634568
rect 127124 634556 127130 634568
rect 132466 634556 132494 634596
rect 155954 634584 155960 634596
rect 156012 634584 156018 634636
rect 165982 634584 165988 634636
rect 166040 634624 166046 634636
rect 177298 634624 177304 634636
rect 166040 634596 177304 634624
rect 166040 634584 166046 634596
rect 177298 634584 177304 634596
rect 177356 634584 177362 634636
rect 183646 634584 183652 634636
rect 183704 634624 183710 634636
rect 211706 634624 211712 634636
rect 183704 634596 211712 634624
rect 183704 634584 183710 634596
rect 211706 634584 211712 634596
rect 211764 634584 211770 634636
rect 221918 634584 221924 634636
rect 221976 634624 221982 634636
rect 232498 634624 232504 634636
rect 221976 634596 232504 634624
rect 221976 634584 221982 634596
rect 232498 634584 232504 634596
rect 232556 634584 232562 634636
rect 238846 634584 238852 634636
rect 238904 634624 238910 634636
rect 268010 634624 268016 634636
rect 238904 634596 268016 634624
rect 238904 634584 238910 634596
rect 268010 634584 268016 634596
rect 268068 634584 268074 634636
rect 277670 634584 277676 634636
rect 277728 634624 277734 634636
rect 289078 634624 289084 634636
rect 277728 634596 289084 634624
rect 277728 634584 277734 634596
rect 289078 634584 289084 634596
rect 289136 634584 289142 634636
rect 306006 634584 306012 634636
rect 306064 634624 306070 634636
rect 316678 634624 316684 634636
rect 306064 634596 316684 634624
rect 306064 634584 306070 634596
rect 316678 634584 316684 634596
rect 316736 634584 316742 634636
rect 323026 634584 323032 634636
rect 323084 634624 323090 634636
rect 352006 634624 352012 634636
rect 323084 634596 352012 634624
rect 323084 634584 323090 634596
rect 352006 634584 352012 634596
rect 352064 634584 352070 634636
rect 361666 634584 361672 634636
rect 361724 634624 361730 634636
rect 373258 634624 373264 634636
rect 361724 634596 373264 634624
rect 361724 634584 361730 634596
rect 373258 634584 373264 634596
rect 373316 634584 373322 634636
rect 379606 634584 379612 634636
rect 379664 634624 379670 634636
rect 408034 634624 408040 634636
rect 379664 634596 408040 634624
rect 379664 634584 379670 634596
rect 408034 634584 408040 634596
rect 408092 634584 408098 634636
rect 417694 634584 417700 634636
rect 417752 634624 417758 634636
rect 428550 634624 428556 634636
rect 417752 634596 428556 634624
rect 417752 634584 417758 634596
rect 428550 634584 428556 634596
rect 428608 634584 428614 634636
rect 434806 634584 434812 634636
rect 434864 634624 434870 634636
rect 463786 634624 463792 634636
rect 434864 634596 463792 634624
rect 434864 634584 434870 634596
rect 463786 634584 463792 634596
rect 463844 634584 463850 634636
rect 473998 634584 474004 634636
rect 474056 634624 474062 634636
rect 485038 634624 485044 634636
rect 474056 634596 485044 634624
rect 474056 634584 474062 634596
rect 485038 634584 485044 634596
rect 485096 634584 485102 634636
rect 501690 634584 501696 634636
rect 501748 634624 501754 634636
rect 512638 634624 512644 634636
rect 501748 634596 512644 634624
rect 501748 634584 501754 634596
rect 512638 634584 512644 634596
rect 512696 634584 512702 634636
rect 518986 634584 518992 634636
rect 519044 634624 519050 634636
rect 547874 634624 547880 634636
rect 519044 634596 547880 634624
rect 519044 634584 519050 634596
rect 547874 634584 547880 634596
rect 547932 634584 547938 634636
rect 127124 634528 132494 634556
rect 127124 634516 127130 634528
rect 137646 634516 137652 634568
rect 137704 634556 137710 634568
rect 148410 634556 148416 634568
rect 137704 634528 148416 634556
rect 137704 634516 137710 634528
rect 148410 634516 148416 634528
rect 148468 634516 148474 634568
rect 193674 634516 193680 634568
rect 193732 634556 193738 634568
rect 204898 634556 204904 634568
rect 193732 634528 204904 634556
rect 193732 634516 193738 634528
rect 204898 634516 204904 634528
rect 204956 634516 204962 634568
rect 249702 634516 249708 634568
rect 249760 634556 249766 634568
rect 260098 634556 260104 634568
rect 249760 634528 260104 634556
rect 249760 634516 249766 634528
rect 260098 634516 260104 634528
rect 260156 634516 260162 634568
rect 333698 634516 333704 634568
rect 333756 634556 333762 634568
rect 344278 634556 344284 634568
rect 333756 634528 344284 634556
rect 333756 634516 333762 634528
rect 344278 634516 344284 634528
rect 344336 634516 344342 634568
rect 390002 634516 390008 634568
rect 390060 634556 390066 634568
rect 400858 634556 400864 634568
rect 390060 634528 400864 634556
rect 390060 634516 390066 634528
rect 400858 634516 400864 634528
rect 400916 634516 400922 634568
rect 445662 634516 445668 634568
rect 445720 634556 445726 634568
rect 456150 634556 456156 634568
rect 445720 634528 456156 634556
rect 445720 634516 445726 634528
rect 456150 634516 456156 634528
rect 456208 634516 456214 634568
rect 529658 634516 529664 634568
rect 529716 634556 529722 634568
rect 540238 634556 540244 634568
rect 529716 634528 540244 634556
rect 529716 634516 529722 634528
rect 540238 634516 540244 634528
rect 540296 634516 540302 634568
rect 36722 634448 36728 634500
rect 36780 634488 36786 634500
rect 557534 634488 557540 634500
rect 36780 634460 557540 634488
rect 36780 634448 36786 634460
rect 557534 634448 557540 634460
rect 557592 634448 557598 634500
rect 16022 632680 16028 632732
rect 16080 632720 16086 632732
rect 547874 632720 547880 632732
rect 16080 632692 547880 632720
rect 16080 632680 16086 632692
rect 547874 632680 547880 632692
rect 547932 632680 547938 632732
rect 25682 632272 25688 632324
rect 25740 632312 25746 632324
rect 71038 632312 71044 632324
rect 25740 632284 71044 632312
rect 25740 632272 25746 632284
rect 71038 632272 71044 632284
rect 71096 632272 71102 632324
rect 212350 632272 212356 632324
rect 212408 632312 212414 632324
rect 232682 632312 232688 632324
rect 212408 632284 232688 632312
rect 212408 632272 212414 632284
rect 232682 632272 232688 632284
rect 232740 632272 232746 632324
rect 408034 632272 408040 632324
rect 408092 632312 408098 632324
rect 428642 632312 428648 632324
rect 408092 632284 428648 632312
rect 408092 632272 408098 632284
rect 428642 632272 428648 632284
rect 428700 632272 428706 632324
rect 492030 632272 492036 632324
rect 492088 632312 492094 632324
rect 512730 632312 512736 632324
rect 492088 632284 512736 632312
rect 492088 632272 492094 632284
rect 512730 632272 512736 632284
rect 512788 632272 512794 632324
rect 36998 632204 37004 632256
rect 37056 632244 37062 632256
rect 53650 632244 53656 632256
rect 37056 632216 53656 632244
rect 37056 632204 37062 632216
rect 53650 632204 53656 632216
rect 53708 632204 53714 632256
rect 148318 632204 148324 632256
rect 148376 632244 148382 632256
rect 165706 632244 165712 632256
rect 148376 632216 165712 632244
rect 148376 632204 148382 632216
rect 165706 632204 165712 632216
rect 165764 632204 165770 632256
rect 175458 632204 175464 632256
rect 175516 632244 175522 632256
rect 193674 632244 193680 632256
rect 175516 632216 193680 632244
rect 175516 632204 175522 632216
rect 193674 632204 193680 632216
rect 193732 632204 193738 632256
rect 203518 632204 203524 632256
rect 203576 632244 203582 632256
rect 221366 632244 221372 632256
rect 203576 632216 221372 632244
rect 203576 632204 203582 632216
rect 221366 632204 221372 632216
rect 221424 632204 221430 632256
rect 260098 632204 260104 632256
rect 260156 632244 260162 632256
rect 277670 632244 277676 632256
rect 260156 632216 277676 632244
rect 260156 632204 260162 632216
rect 277670 632204 277676 632216
rect 277728 632204 277734 632256
rect 287514 632204 287520 632256
rect 287572 632244 287578 632256
rect 305362 632244 305368 632256
rect 287572 632216 305368 632244
rect 287572 632204 287578 632216
rect 305362 632204 305368 632216
rect 305420 632204 305426 632256
rect 315482 632204 315488 632256
rect 315540 632244 315546 632256
rect 333698 632244 333704 632256
rect 315540 632216 333704 632244
rect 315540 632204 315546 632216
rect 333698 632204 333704 632216
rect 333756 632204 333762 632256
rect 345658 632204 345664 632256
rect 345716 632244 345722 632256
rect 361666 632244 361672 632256
rect 345716 632216 361672 632244
rect 345716 632204 345722 632216
rect 361666 632204 361672 632216
rect 361724 632204 361730 632256
rect 371510 632204 371516 632256
rect 371568 632244 371574 632256
rect 389358 632244 389364 632256
rect 371568 632216 389364 632244
rect 371568 632204 371574 632216
rect 389358 632204 389364 632216
rect 389416 632204 389422 632256
rect 399478 632204 399484 632256
rect 399536 632244 399542 632256
rect 417694 632244 417700 632256
rect 399536 632216 417700 632244
rect 399536 632204 399542 632216
rect 417694 632204 417700 632216
rect 417752 632204 417758 632256
rect 456150 632204 456156 632256
rect 456208 632244 456214 632256
rect 473354 632244 473360 632256
rect 456208 632216 473360 632244
rect 456208 632204 456214 632216
rect 473354 632204 473360 632216
rect 473412 632204 473418 632256
rect 483474 632204 483480 632256
rect 483532 632244 483538 632256
rect 501690 632244 501696 632256
rect 483532 632216 501696 632244
rect 483532 632204 483538 632216
rect 501690 632204 501696 632216
rect 501748 632204 501754 632256
rect 36906 632136 36912 632188
rect 36964 632176 36970 632188
rect 63310 632176 63316 632188
rect 36964 632148 63316 632176
rect 36964 632136 36970 632148
rect 63310 632136 63316 632148
rect 63368 632136 63374 632188
rect 64322 632136 64328 632188
rect 64380 632176 64386 632188
rect 81434 632176 81440 632188
rect 64380 632148 81440 632176
rect 64380 632136 64386 632148
rect 81434 632136 81440 632148
rect 81492 632136 81498 632188
rect 91462 632136 91468 632188
rect 91520 632176 91526 632188
rect 109678 632176 109684 632188
rect 91520 632148 109684 632176
rect 91520 632136 91526 632148
rect 109678 632136 109684 632148
rect 109736 632136 109742 632188
rect 119430 632136 119436 632188
rect 119488 632176 119494 632188
rect 137646 632176 137652 632188
rect 119488 632148 137652 632176
rect 119488 632136 119494 632148
rect 137646 632136 137652 632148
rect 137704 632136 137710 632188
rect 156322 632136 156328 632188
rect 156380 632176 156386 632188
rect 178678 632176 178684 632188
rect 156380 632148 178684 632176
rect 156380 632136 156386 632148
rect 178678 632136 178684 632148
rect 178736 632136 178742 632188
rect 232590 632136 232596 632188
rect 232648 632176 232654 632188
rect 249702 632176 249708 632188
rect 232648 632148 249708 632176
rect 232648 632136 232654 632148
rect 249702 632136 249708 632148
rect 249760 632136 249766 632188
rect 268010 632136 268016 632188
rect 268068 632176 268074 632188
rect 287698 632176 287704 632188
rect 268068 632148 287704 632176
rect 268068 632136 268074 632148
rect 287698 632136 287704 632148
rect 287756 632136 287762 632188
rect 296346 632136 296352 632188
rect 296404 632176 296410 632188
rect 316770 632176 316776 632188
rect 296404 632148 316776 632176
rect 296404 632136 296410 632148
rect 316770 632136 316776 632148
rect 316828 632136 316834 632188
rect 352006 632136 352012 632188
rect 352064 632176 352070 632188
rect 374638 632176 374644 632188
rect 352064 632148 374644 632176
rect 352064 632136 352070 632148
rect 374638 632136 374644 632148
rect 374696 632136 374702 632188
rect 428458 632136 428464 632188
rect 428516 632176 428522 632188
rect 445662 632176 445668 632188
rect 428516 632148 445668 632176
rect 428516 632136 428522 632148
rect 445662 632136 445668 632148
rect 445720 632136 445726 632188
rect 464338 632136 464344 632188
rect 464396 632176 464402 632188
rect 483658 632176 483664 632188
rect 464396 632148 483664 632176
rect 464396 632136 464402 632148
rect 483658 632136 483664 632148
rect 483716 632136 483722 632188
rect 511442 632136 511448 632188
rect 511500 632176 511506 632188
rect 529658 632176 529664 632188
rect 511500 632148 529664 632176
rect 511500 632136 511506 632148
rect 529658 632136 529664 632148
rect 529716 632136 529722 632188
rect 542998 632136 543004 632188
rect 543056 632176 543062 632188
rect 557534 632176 557540 632188
rect 543056 632148 557540 632176
rect 543056 632136 543062 632148
rect 557534 632136 557540 632148
rect 557592 632136 557598 632188
rect 3142 632068 3148 632120
rect 3200 632108 3206 632120
rect 6178 632108 6184 632120
rect 3200 632080 6184 632108
rect 3200 632068 3206 632080
rect 6178 632068 6184 632080
rect 6236 632068 6242 632120
rect 69658 632068 69664 632120
rect 69716 632108 69722 632120
rect 91094 632108 91100 632120
rect 69716 632080 91100 632108
rect 69716 632068 69722 632080
rect 91094 632068 91100 632080
rect 91152 632068 91158 632120
rect 95878 632068 95884 632120
rect 95936 632108 95942 632120
rect 119338 632108 119344 632120
rect 95936 632080 119344 632108
rect 95936 632068 95942 632080
rect 119338 632068 119344 632080
rect 119396 632068 119402 632120
rect 120718 632068 120724 632120
rect 120776 632108 120782 632120
rect 147306 632108 147312 632120
rect 120776 632080 147312 632108
rect 120776 632068 120782 632080
rect 147306 632068 147312 632080
rect 147364 632068 147370 632120
rect 148410 632068 148416 632120
rect 148468 632108 148474 632120
rect 175366 632108 175372 632120
rect 148468 632080 175372 632108
rect 148468 632068 148474 632080
rect 175366 632068 175372 632080
rect 175424 632068 175430 632120
rect 177298 632068 177304 632120
rect 177356 632108 177362 632120
rect 203334 632108 203340 632120
rect 177356 632080 203340 632108
rect 177356 632068 177362 632080
rect 203334 632068 203340 632080
rect 203392 632068 203398 632120
rect 204898 632068 204904 632120
rect 204956 632108 204962 632120
rect 231026 632108 231032 632120
rect 204956 632080 231032 632108
rect 204956 632068 204962 632080
rect 231026 632068 231032 632080
rect 231084 632068 231090 632120
rect 232498 632068 232504 632120
rect 232556 632108 232562 632120
rect 259362 632108 259368 632120
rect 232556 632080 259368 632108
rect 232556 632068 232562 632080
rect 259362 632068 259368 632080
rect 259420 632068 259426 632120
rect 260190 632068 260196 632120
rect 260248 632108 260254 632120
rect 287330 632108 287336 632120
rect 260248 632080 287336 632108
rect 260248 632068 260254 632080
rect 287330 632068 287336 632080
rect 287388 632068 287394 632120
rect 289078 632068 289084 632120
rect 289136 632108 289142 632120
rect 315022 632108 315028 632120
rect 289136 632080 315028 632108
rect 289136 632068 289142 632080
rect 315022 632068 315028 632080
rect 315080 632068 315086 632120
rect 316678 632068 316684 632120
rect 316736 632108 316742 632120
rect 343358 632108 343364 632120
rect 316736 632080 343364 632108
rect 316736 632068 316742 632080
rect 343358 632068 343364 632080
rect 343416 632068 343422 632120
rect 344278 632068 344284 632120
rect 344336 632108 344342 632120
rect 371326 632108 371332 632120
rect 344336 632080 371332 632108
rect 344336 632068 344342 632080
rect 371326 632068 371332 632080
rect 371384 632068 371390 632120
rect 373258 632068 373264 632120
rect 373316 632108 373322 632120
rect 399018 632108 399024 632120
rect 373316 632080 399024 632108
rect 373316 632068 373322 632080
rect 399018 632068 399024 632080
rect 399076 632068 399082 632120
rect 400858 632068 400864 632120
rect 400916 632108 400922 632120
rect 427354 632108 427360 632120
rect 400916 632080 427360 632108
rect 400916 632068 400922 632080
rect 427354 632068 427360 632080
rect 427412 632068 427418 632120
rect 428550 632068 428556 632120
rect 428608 632108 428614 632120
rect 455322 632108 455328 632120
rect 428608 632080 455328 632108
rect 428608 632068 428614 632080
rect 455322 632068 455328 632080
rect 455380 632068 455386 632120
rect 456058 632068 456064 632120
rect 456116 632108 456122 632120
rect 483014 632108 483020 632120
rect 456116 632080 483020 632108
rect 456116 632068 456122 632080
rect 483014 632068 483020 632080
rect 483072 632068 483078 632120
rect 485038 632068 485044 632120
rect 485096 632108 485102 632120
rect 511350 632108 511356 632120
rect 485096 632080 511356 632108
rect 485096 632068 485102 632080
rect 511350 632068 511356 632080
rect 511408 632068 511414 632120
rect 512638 632068 512644 632120
rect 512696 632108 512702 632120
rect 539318 632108 539324 632120
rect 512696 632080 539324 632108
rect 512696 632068 512702 632080
rect 539318 632068 539324 632080
rect 539376 632068 539382 632120
rect 540238 632068 540244 632120
rect 540296 632108 540302 632120
rect 567194 632108 567200 632120
rect 540296 632080 567200 632108
rect 540296 632068 540302 632080
rect 567194 632068 567200 632080
rect 567252 632068 567258 632120
rect 37918 629892 37924 629944
rect 37976 629932 37982 629944
rect 545758 629932 545764 629944
rect 37976 629904 545764 629932
rect 37976 629892 37982 629904
rect 545758 629892 545764 629904
rect 545816 629892 545822 629944
rect 35618 629280 35624 629332
rect 35676 629320 35682 629332
rect 36722 629320 36728 629332
rect 35676 629292 36728 629320
rect 35676 629280 35682 629292
rect 36722 629280 36728 629292
rect 36780 629280 36786 629332
rect 567930 616836 567936 616888
rect 567988 616876 567994 616888
rect 580166 616876 580172 616888
rect 567988 616848 580172 616876
rect 567988 616836 567994 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 63586 612756 63592 612808
rect 63644 612796 63650 612808
rect 64322 612796 64328 612808
rect 63644 612768 64328 612796
rect 63644 612756 63650 612768
rect 64322 612756 64328 612768
rect 64380 612756 64386 612808
rect 455690 612756 455696 612808
rect 455748 612796 455754 612808
rect 456150 612796 456156 612808
rect 455748 612768 456156 612796
rect 455748 612756 455754 612768
rect 456150 612756 456156 612768
rect 456208 612756 456214 612808
rect 316770 612008 316776 612060
rect 316828 612048 316834 612060
rect 323670 612048 323676 612060
rect 316828 612020 323676 612048
rect 316828 612008 316834 612020
rect 323670 612008 323676 612020
rect 323728 612008 323734 612060
rect 428642 612008 428648 612060
rect 428700 612048 428706 612060
rect 435726 612048 435732 612060
rect 428700 612020 435732 612048
rect 428700 612008 428706 612020
rect 435726 612008 435732 612020
rect 435784 612008 435790 612060
rect 232682 611940 232688 611992
rect 232740 611980 232746 611992
rect 239766 611980 239772 611992
rect 232740 611952 239772 611980
rect 232740 611940 232746 611952
rect 239766 611940 239772 611952
rect 239824 611940 239830 611992
rect 287698 611872 287704 611924
rect 287756 611912 287762 611924
rect 295702 611912 295708 611924
rect 287756 611884 295708 611912
rect 287756 611872 287762 611884
rect 295702 611872 295708 611884
rect 295760 611872 295766 611924
rect 483658 611736 483664 611788
rect 483716 611776 483722 611788
rect 491662 611776 491668 611788
rect 483716 611748 491668 611776
rect 483716 611736 483722 611748
rect 491662 611736 491668 611748
rect 491720 611736 491726 611788
rect 512730 611736 512736 611788
rect 512788 611776 512794 611788
rect 519630 611776 519636 611788
rect 512788 611748 519636 611776
rect 512788 611736 512794 611748
rect 519630 611736 519636 611748
rect 519688 611736 519694 611788
rect 13722 611260 13728 611312
rect 13780 611300 13786 611312
rect 66254 611300 66260 611312
rect 13780 611272 66260 611300
rect 13780 611260 13786 611272
rect 66254 611260 66260 611272
rect 66312 611260 66318 611312
rect 70302 611260 70308 611312
rect 70360 611300 70366 611312
rect 121454 611300 121460 611312
rect 70360 611272 121460 611300
rect 70360 611260 70366 611272
rect 121454 611260 121460 611272
rect 121512 611260 121518 611312
rect 126882 611260 126888 611312
rect 126940 611300 126946 611312
rect 178034 611300 178040 611312
rect 126940 611272 178040 611300
rect 126940 611260 126946 611272
rect 178034 611260 178040 611272
rect 178092 611260 178098 611312
rect 209682 611260 209688 611312
rect 209740 611300 209746 611312
rect 262214 611300 262220 611312
rect 209740 611272 262220 611300
rect 209740 611260 209746 611272
rect 262214 611260 262220 611272
rect 262272 611260 262278 611312
rect 266262 611260 266268 611312
rect 266320 611300 266326 611312
rect 317414 611300 317420 611312
rect 266320 611272 317420 611300
rect 266320 611260 266326 611272
rect 317414 611260 317420 611272
rect 317472 611260 317478 611312
rect 322842 611260 322848 611312
rect 322900 611300 322906 611312
rect 373994 611300 374000 611312
rect 322900 611272 374000 611300
rect 322900 611260 322906 611272
rect 373994 611260 374000 611272
rect 374052 611260 374058 611312
rect 405642 611260 405648 611312
rect 405700 611300 405706 611312
rect 458174 611300 458180 611312
rect 405700 611272 458180 611300
rect 405700 611260 405706 611272
rect 458174 611260 458180 611272
rect 458232 611260 458238 611312
rect 489822 611260 489828 611312
rect 489880 611300 489886 611312
rect 542354 611300 542360 611312
rect 489880 611272 542360 611300
rect 489880 611260 489886 611272
rect 542354 611260 542360 611272
rect 542412 611260 542418 611312
rect 35618 611192 35624 611244
rect 35676 611232 35682 611244
rect 36998 611232 37004 611244
rect 35676 611204 37004 611232
rect 35676 611192 35682 611204
rect 36998 611192 37004 611204
rect 37056 611192 37062 611244
rect 42702 611192 42708 611244
rect 42760 611232 42766 611244
rect 93854 611232 93860 611244
rect 42760 611204 93860 611232
rect 42760 611192 42766 611204
rect 93854 611192 93860 611204
rect 93912 611192 93918 611244
rect 97902 611192 97908 611244
rect 97960 611232 97966 611244
rect 149054 611232 149060 611244
rect 97960 611204 149060 611232
rect 97960 611192 97966 611204
rect 149054 611192 149060 611204
rect 149112 611192 149118 611244
rect 154482 611192 154488 611244
rect 154540 611232 154546 611244
rect 205634 611232 205640 611244
rect 154540 611204 205640 611232
rect 154540 611192 154546 611204
rect 205634 611192 205640 611204
rect 205692 611192 205698 611244
rect 231670 611192 231676 611244
rect 231728 611232 231734 611244
rect 232590 611232 232596 611244
rect 231728 611204 232596 611232
rect 231728 611192 231734 611204
rect 232590 611192 232596 611204
rect 232648 611192 232654 611244
rect 238662 611192 238668 611244
rect 238720 611232 238726 611244
rect 289814 611232 289820 611244
rect 238720 611204 289820 611232
rect 238720 611192 238726 611204
rect 289814 611192 289820 611204
rect 289872 611192 289878 611244
rect 293862 611192 293868 611244
rect 293920 611232 293926 611244
rect 345014 611232 345020 611244
rect 293920 611204 345020 611232
rect 293920 611192 293926 611204
rect 345014 611192 345020 611204
rect 345072 611192 345078 611244
rect 350442 611192 350448 611244
rect 350500 611232 350506 611244
rect 401594 611232 401600 611244
rect 350500 611204 401600 611232
rect 350500 611192 350506 611204
rect 401594 611192 401600 611204
rect 401652 611192 401658 611244
rect 462222 611192 462228 611244
rect 462280 611232 462286 611244
rect 513374 611232 513380 611244
rect 462280 611204 513380 611232
rect 462280 611192 462286 611204
rect 513374 611192 513380 611204
rect 513432 611192 513438 611244
rect 518802 611192 518808 611244
rect 518860 611232 518866 611244
rect 569954 611232 569960 611244
rect 518860 611204 569960 611232
rect 518860 611192 518866 611204
rect 569954 611192 569960 611204
rect 570012 611192 570018 611244
rect 182082 611124 182088 611176
rect 182140 611164 182146 611176
rect 233234 611164 233240 611176
rect 182140 611136 233240 611164
rect 182140 611124 182146 611136
rect 233234 611124 233240 611136
rect 233292 611124 233298 611176
rect 378042 611124 378048 611176
rect 378100 611164 378106 611176
rect 429194 611164 429200 611176
rect 378100 611136 429200 611164
rect 378100 611124 378106 611136
rect 429194 611124 429200 611136
rect 429252 611124 429258 611176
rect 434622 611124 434628 611176
rect 434680 611164 434686 611176
rect 485774 611164 485780 611176
rect 434680 611136 485780 611164
rect 434680 611124 434686 611136
rect 485774 611124 485780 611136
rect 485832 611124 485838 611176
rect 72050 608580 72056 608592
rect 64846 608552 72056 608580
rect 15194 608472 15200 608524
rect 15252 608512 15258 608524
rect 43990 608512 43996 608524
rect 15252 608484 43996 608512
rect 15252 608472 15258 608484
rect 43990 608472 43996 608484
rect 44048 608472 44054 608524
rect 25682 608404 25688 608456
rect 25740 608444 25746 608456
rect 36906 608444 36912 608456
rect 25740 608416 36912 608444
rect 25740 608404 25746 608416
rect 36906 608404 36912 608416
rect 36964 608404 36970 608456
rect 42886 608404 42892 608456
rect 42944 608444 42950 608456
rect 64846 608444 64874 608552
rect 72050 608540 72056 608552
rect 72108 608540 72114 608592
rect 178678 608540 178684 608592
rect 178736 608580 178742 608592
rect 184014 608580 184020 608592
rect 178736 608552 184020 608580
rect 178736 608540 178742 608552
rect 184014 608540 184020 608552
rect 184072 608540 184078 608592
rect 343358 608540 343364 608592
rect 343416 608580 343422 608592
rect 345658 608580 345664 608592
rect 343416 608552 345664 608580
rect 343416 608540 343422 608552
rect 345658 608540 345664 608552
rect 345716 608540 345722 608592
rect 374638 608540 374644 608592
rect 374696 608580 374702 608592
rect 379698 608580 379704 608592
rect 374696 608552 379704 608580
rect 374696 608540 374702 608552
rect 379698 608540 379704 608552
rect 379756 608540 379762 608592
rect 539318 608540 539324 608592
rect 539376 608580 539382 608592
rect 542998 608580 543004 608592
rect 539376 608552 543004 608580
rect 539376 608540 539382 608552
rect 542998 608540 543004 608552
rect 543056 608540 543062 608592
rect 66898 608472 66904 608524
rect 66956 608512 66962 608524
rect 567194 608512 567200 608524
rect 66956 608484 567200 608512
rect 66956 608472 66962 608484
rect 567194 608472 567200 608484
rect 567252 608472 567258 608524
rect 42944 608416 64874 608444
rect 42944 608404 42950 608416
rect 71866 608404 71872 608456
rect 71924 608444 71930 608456
rect 100018 608444 100024 608456
rect 71924 608416 100024 608444
rect 71924 608404 71930 608416
rect 100018 608404 100024 608416
rect 100076 608404 100082 608456
rect 127986 608444 127992 608456
rect 103486 608416 127992 608444
rect 53650 608336 53656 608388
rect 53708 608376 53714 608388
rect 69658 608376 69664 608388
rect 53708 608348 69664 608376
rect 53708 608336 53714 608348
rect 69658 608336 69664 608348
rect 69716 608336 69722 608388
rect 81986 608336 81992 608388
rect 82044 608376 82050 608388
rect 95878 608376 95884 608388
rect 82044 608348 95884 608376
rect 82044 608336 82050 608348
rect 95878 608336 95884 608348
rect 95936 608336 95942 608388
rect 99466 608336 99472 608388
rect 99524 608376 99530 608388
rect 103486 608376 103514 608416
rect 127986 608404 127992 608416
rect 128044 608404 128050 608456
rect 156046 608444 156052 608456
rect 132466 608416 156052 608444
rect 99524 608348 103514 608376
rect 99524 608336 99530 608348
rect 109678 608336 109684 608388
rect 109736 608376 109742 608388
rect 120718 608376 120724 608388
rect 109736 608348 120724 608376
rect 109736 608336 109742 608348
rect 120718 608336 120724 608348
rect 120776 608336 120782 608388
rect 127066 608336 127072 608388
rect 127124 608376 127130 608388
rect 132466 608376 132494 608416
rect 156046 608404 156052 608416
rect 156104 608404 156110 608456
rect 165982 608404 165988 608456
rect 166040 608444 166046 608456
rect 177298 608444 177304 608456
rect 166040 608416 177304 608444
rect 166040 608404 166046 608416
rect 177298 608404 177304 608416
rect 177356 608404 177362 608456
rect 183646 608404 183652 608456
rect 183704 608444 183710 608456
rect 211706 608444 211712 608456
rect 183704 608416 211712 608444
rect 183704 608404 183710 608416
rect 211706 608404 211712 608416
rect 211764 608404 211770 608456
rect 222010 608404 222016 608456
rect 222068 608444 222074 608456
rect 232498 608444 232504 608456
rect 222068 608416 232504 608444
rect 222068 608404 222074 608416
rect 232498 608404 232504 608416
rect 232556 608404 232562 608456
rect 238846 608404 238852 608456
rect 238904 608444 238910 608456
rect 268010 608444 268016 608456
rect 238904 608416 268016 608444
rect 238904 608404 238910 608416
rect 268010 608404 268016 608416
rect 268068 608404 268074 608456
rect 277670 608404 277676 608456
rect 277728 608444 277734 608456
rect 289078 608444 289084 608456
rect 277728 608416 289084 608444
rect 277728 608404 277734 608416
rect 289078 608404 289084 608416
rect 289136 608404 289142 608456
rect 306006 608404 306012 608456
rect 306064 608444 306070 608456
rect 316678 608444 316684 608456
rect 306064 608416 316684 608444
rect 306064 608404 306070 608416
rect 316678 608404 316684 608416
rect 316736 608404 316742 608456
rect 323026 608404 323032 608456
rect 323084 608444 323090 608456
rect 352006 608444 352012 608456
rect 323084 608416 352012 608444
rect 323084 608404 323090 608416
rect 352006 608404 352012 608416
rect 352064 608404 352070 608456
rect 361666 608404 361672 608456
rect 361724 608444 361730 608456
rect 373258 608444 373264 608456
rect 361724 608416 373264 608444
rect 361724 608404 361730 608416
rect 373258 608404 373264 608416
rect 373316 608404 373322 608456
rect 379606 608404 379612 608456
rect 379664 608444 379670 608456
rect 408034 608444 408040 608456
rect 379664 608416 408040 608444
rect 379664 608404 379670 608416
rect 408034 608404 408040 608416
rect 408092 608404 408098 608456
rect 417694 608404 417700 608456
rect 417752 608444 417758 608456
rect 428550 608444 428556 608456
rect 417752 608416 428556 608444
rect 417752 608404 417758 608416
rect 428550 608404 428556 608416
rect 428608 608404 428614 608456
rect 434806 608404 434812 608456
rect 434864 608444 434870 608456
rect 463694 608444 463700 608456
rect 434864 608416 463700 608444
rect 434864 608404 434870 608416
rect 463694 608404 463700 608416
rect 463752 608404 463758 608456
rect 473998 608404 474004 608456
rect 474056 608444 474062 608456
rect 485038 608444 485044 608456
rect 474056 608416 485044 608444
rect 474056 608404 474062 608416
rect 485038 608404 485044 608416
rect 485096 608404 485102 608456
rect 501690 608404 501696 608456
rect 501748 608444 501754 608456
rect 512638 608444 512644 608456
rect 501748 608416 512644 608444
rect 501748 608404 501754 608416
rect 512638 608404 512644 608416
rect 512696 608404 512702 608456
rect 518986 608404 518992 608456
rect 519044 608444 519050 608456
rect 547874 608444 547880 608456
rect 519044 608416 547880 608444
rect 519044 608404 519050 608416
rect 547874 608404 547880 608416
rect 547932 608404 547938 608456
rect 127124 608348 132494 608376
rect 127124 608336 127130 608348
rect 137646 608336 137652 608388
rect 137704 608376 137710 608388
rect 148410 608376 148416 608388
rect 137704 608348 148416 608376
rect 137704 608336 137710 608348
rect 148410 608336 148416 608348
rect 148468 608336 148474 608388
rect 193674 608336 193680 608388
rect 193732 608376 193738 608388
rect 204898 608376 204904 608388
rect 193732 608348 204904 608376
rect 193732 608336 193738 608348
rect 204898 608336 204904 608348
rect 204956 608336 204962 608388
rect 249702 608336 249708 608388
rect 249760 608376 249766 608388
rect 260190 608376 260196 608388
rect 249760 608348 260196 608376
rect 249760 608336 249766 608348
rect 260190 608336 260196 608348
rect 260248 608336 260254 608388
rect 333698 608336 333704 608388
rect 333756 608376 333762 608388
rect 344278 608376 344284 608388
rect 333756 608348 344284 608376
rect 333756 608336 333762 608348
rect 344278 608336 344284 608348
rect 344336 608336 344342 608388
rect 390002 608336 390008 608388
rect 390060 608376 390066 608388
rect 400858 608376 400864 608388
rect 390060 608348 400864 608376
rect 390060 608336 390066 608348
rect 400858 608336 400864 608348
rect 400916 608336 400922 608388
rect 445662 608336 445668 608388
rect 445720 608376 445726 608388
rect 456058 608376 456064 608388
rect 445720 608348 456064 608376
rect 445720 608336 445726 608348
rect 456058 608336 456064 608348
rect 456116 608336 456122 608388
rect 529658 608336 529664 608388
rect 529716 608376 529722 608388
rect 540238 608376 540244 608388
rect 529716 608348 540244 608376
rect 529716 608336 529722 608348
rect 540238 608336 540244 608348
rect 540296 608336 540302 608388
rect 36814 608268 36820 608320
rect 36872 608308 36878 608320
rect 557534 608308 557540 608320
rect 36872 608280 557540 608308
rect 36872 608268 36878 608280
rect 557534 608268 557540 608280
rect 557592 608268 557598 608320
rect 15286 605072 15292 605124
rect 15344 605112 15350 605124
rect 547874 605112 547880 605124
rect 15344 605084 547880 605112
rect 15344 605072 15350 605084
rect 547874 605072 547880 605084
rect 547932 605072 547938 605124
rect 25682 604732 25688 604784
rect 25740 604772 25746 604784
rect 261478 604772 261484 604784
rect 25740 604744 261484 604772
rect 25740 604732 25746 604744
rect 261478 604732 261484 604744
rect 261536 604732 261542 604784
rect 119430 604664 119436 604716
rect 119488 604704 119494 604716
rect 137646 604704 137652 604716
rect 119488 604676 137652 604704
rect 119488 604664 119494 604676
rect 137646 604664 137652 604676
rect 137704 604664 137710 604716
rect 148318 604664 148324 604716
rect 148376 604704 148382 604716
rect 165706 604704 165712 604716
rect 148376 604676 165712 604704
rect 148376 604664 148382 604676
rect 165706 604664 165712 604676
rect 165764 604664 165770 604716
rect 175458 604664 175464 604716
rect 175516 604704 175522 604716
rect 193674 604704 193680 604716
rect 175516 604676 193680 604704
rect 175516 604664 175522 604676
rect 193674 604664 193680 604676
rect 193732 604664 193738 604716
rect 203518 604664 203524 604716
rect 203576 604704 203582 604716
rect 221366 604704 221372 604716
rect 203576 604676 221372 604704
rect 203576 604664 203582 604676
rect 221366 604664 221372 604676
rect 221424 604664 221430 604716
rect 408034 604664 408040 604716
rect 408092 604704 408098 604716
rect 428642 604704 428648 604716
rect 408092 604676 428648 604704
rect 408092 604664 408098 604676
rect 428642 604664 428648 604676
rect 428700 604664 428706 604716
rect 492030 604664 492036 604716
rect 492088 604704 492094 604716
rect 512730 604704 512736 604716
rect 492088 604676 512736 604704
rect 492088 604664 492094 604676
rect 512730 604664 512736 604676
rect 512788 604664 512794 604716
rect 36998 604596 37004 604648
rect 37056 604636 37062 604648
rect 53650 604636 53656 604648
rect 37056 604608 53656 604636
rect 37056 604596 37062 604608
rect 53650 604596 53656 604608
rect 53708 604596 53714 604648
rect 64322 604596 64328 604648
rect 64380 604636 64386 604648
rect 81434 604636 81440 604648
rect 64380 604608 81440 604636
rect 64380 604596 64386 604608
rect 81434 604596 81440 604608
rect 81492 604596 81498 604648
rect 91462 604596 91468 604648
rect 91520 604636 91526 604648
rect 109678 604636 109684 604648
rect 91520 604608 109684 604636
rect 91520 604596 91526 604608
rect 109678 604596 109684 604608
rect 109736 604596 109742 604648
rect 127986 604596 127992 604648
rect 128044 604636 128050 604648
rect 148502 604636 148508 604648
rect 128044 604608 148508 604636
rect 128044 604596 128050 604608
rect 148502 604596 148508 604608
rect 148560 604596 148566 604648
rect 156322 604596 156328 604648
rect 156380 604636 156386 604648
rect 178678 604636 178684 604648
rect 156380 604608 178684 604636
rect 156380 604596 156386 604608
rect 178678 604596 178684 604608
rect 178736 604596 178742 604648
rect 232498 604596 232504 604648
rect 232556 604636 232562 604648
rect 249702 604636 249708 604648
rect 232556 604608 249708 604636
rect 232556 604596 232562 604608
rect 249702 604596 249708 604608
rect 249760 604596 249766 604648
rect 260190 604596 260196 604648
rect 260248 604636 260254 604648
rect 277670 604636 277676 604648
rect 260248 604608 277676 604636
rect 260248 604596 260254 604608
rect 277670 604596 277676 604608
rect 277728 604596 277734 604648
rect 287514 604596 287520 604648
rect 287572 604636 287578 604648
rect 305362 604636 305368 604648
rect 287572 604608 305368 604636
rect 287572 604596 287578 604608
rect 305362 604596 305368 604608
rect 305420 604596 305426 604648
rect 315482 604596 315488 604648
rect 315540 604636 315546 604648
rect 333698 604636 333704 604648
rect 315540 604608 333704 604636
rect 315540 604596 315546 604608
rect 333698 604596 333704 604608
rect 333756 604596 333762 604648
rect 345658 604596 345664 604648
rect 345716 604636 345722 604648
rect 361666 604636 361672 604648
rect 345716 604608 361672 604636
rect 345716 604596 345722 604608
rect 361666 604596 361672 604608
rect 361724 604596 361730 604648
rect 371510 604596 371516 604648
rect 371568 604636 371574 604648
rect 389358 604636 389364 604648
rect 371568 604608 389364 604636
rect 371568 604596 371574 604608
rect 389358 604596 389364 604608
rect 389416 604596 389422 604648
rect 399478 604596 399484 604648
rect 399536 604636 399542 604648
rect 417694 604636 417700 604648
rect 399536 604608 417700 604636
rect 399536 604596 399542 604608
rect 417694 604596 417700 604608
rect 417752 604596 417758 604648
rect 456058 604596 456064 604648
rect 456116 604636 456122 604648
rect 473354 604636 473360 604648
rect 456116 604608 473360 604636
rect 456116 604596 456122 604608
rect 473354 604596 473360 604608
rect 473412 604596 473418 604648
rect 483474 604596 483480 604648
rect 483532 604636 483538 604648
rect 501690 604636 501696 604648
rect 483532 604608 501696 604636
rect 483532 604596 483538 604608
rect 501690 604596 501696 604608
rect 501748 604596 501754 604648
rect 36906 604528 36912 604580
rect 36964 604568 36970 604580
rect 63310 604568 63316 604580
rect 36964 604540 63316 604568
rect 36964 604528 36970 604540
rect 63310 604528 63316 604540
rect 63368 604528 63374 604580
rect 66898 604528 66904 604580
rect 66956 604568 66962 604580
rect 91094 604568 91100 604580
rect 66956 604540 91100 604568
rect 66956 604528 66962 604540
rect 91094 604528 91100 604540
rect 91152 604528 91158 604580
rect 94498 604528 94504 604580
rect 94556 604568 94562 604580
rect 119338 604568 119344 604580
rect 94556 604540 119344 604568
rect 94556 604528 94562 604540
rect 119338 604528 119344 604540
rect 119396 604528 119402 604580
rect 120718 604528 120724 604580
rect 120776 604568 120782 604580
rect 147306 604568 147312 604580
rect 120776 604540 147312 604568
rect 120776 604528 120782 604540
rect 147306 604528 147312 604540
rect 147364 604528 147370 604580
rect 148410 604528 148416 604580
rect 148468 604568 148474 604580
rect 175366 604568 175372 604580
rect 148468 604540 175372 604568
rect 148468 604528 148474 604540
rect 175366 604528 175372 604540
rect 175424 604528 175430 604580
rect 177298 604528 177304 604580
rect 177356 604568 177362 604580
rect 203334 604568 203340 604580
rect 177356 604540 203340 604568
rect 177356 604528 177362 604540
rect 203334 604528 203340 604540
rect 203392 604528 203398 604580
rect 204898 604528 204904 604580
rect 204956 604568 204962 604580
rect 231026 604568 231032 604580
rect 204956 604540 231032 604568
rect 204956 604528 204962 604540
rect 231026 604528 231032 604540
rect 231084 604528 231090 604580
rect 232590 604528 232596 604580
rect 232648 604568 232654 604580
rect 259362 604568 259368 604580
rect 232648 604540 259368 604568
rect 232648 604528 232654 604540
rect 259362 604528 259368 604540
rect 259420 604528 259426 604580
rect 268010 604528 268016 604580
rect 268068 604568 268074 604580
rect 287698 604568 287704 604580
rect 268068 604540 287704 604568
rect 268068 604528 268074 604540
rect 287698 604528 287704 604540
rect 287756 604528 287762 604580
rect 296346 604528 296352 604580
rect 296404 604568 296410 604580
rect 316770 604568 316776 604580
rect 296404 604540 316776 604568
rect 296404 604528 296410 604540
rect 316770 604528 316776 604540
rect 316828 604528 316834 604580
rect 352006 604528 352012 604580
rect 352064 604568 352070 604580
rect 374638 604568 374644 604580
rect 352064 604540 374644 604568
rect 352064 604528 352070 604540
rect 374638 604528 374644 604540
rect 374696 604528 374702 604580
rect 428550 604528 428556 604580
rect 428608 604568 428614 604580
rect 445662 604568 445668 604580
rect 428608 604540 445668 604568
rect 428608 604528 428614 604540
rect 445662 604528 445668 604540
rect 445720 604528 445726 604580
rect 464338 604528 464344 604580
rect 464396 604568 464402 604580
rect 483658 604568 483664 604580
rect 464396 604540 483664 604568
rect 464396 604528 464402 604540
rect 483658 604528 483664 604540
rect 483716 604528 483722 604580
rect 511442 604528 511448 604580
rect 511500 604568 511506 604580
rect 529658 604568 529664 604580
rect 511500 604540 529664 604568
rect 511500 604528 511506 604540
rect 529658 604528 529664 604540
rect 529716 604528 529722 604580
rect 542998 604528 543004 604580
rect 543056 604568 543062 604580
rect 557534 604568 557540 604580
rect 543056 604540 557540 604568
rect 543056 604528 543062 604540
rect 557534 604528 557540 604540
rect 557592 604528 557598 604580
rect 212350 604460 212356 604512
rect 212408 604500 212414 604512
rect 232682 604500 232688 604512
rect 212408 604472 232688 604500
rect 212408 604460 212414 604472
rect 232682 604460 232688 604472
rect 232740 604460 232746 604512
rect 260098 604460 260104 604512
rect 260156 604500 260162 604512
rect 287330 604500 287336 604512
rect 260156 604472 287336 604500
rect 260156 604460 260162 604472
rect 287330 604460 287336 604472
rect 287388 604460 287394 604512
rect 289078 604460 289084 604512
rect 289136 604500 289142 604512
rect 315022 604500 315028 604512
rect 289136 604472 315028 604500
rect 289136 604460 289142 604472
rect 315022 604460 315028 604472
rect 315080 604460 315086 604512
rect 316678 604460 316684 604512
rect 316736 604500 316742 604512
rect 343358 604500 343364 604512
rect 316736 604472 343364 604500
rect 316736 604460 316742 604472
rect 343358 604460 343364 604472
rect 343416 604460 343422 604512
rect 344278 604460 344284 604512
rect 344336 604500 344342 604512
rect 371326 604500 371332 604512
rect 344336 604472 371332 604500
rect 344336 604460 344342 604472
rect 371326 604460 371332 604472
rect 371384 604460 371390 604512
rect 373258 604460 373264 604512
rect 373316 604500 373322 604512
rect 399018 604500 399024 604512
rect 373316 604472 399024 604500
rect 373316 604460 373322 604472
rect 399018 604460 399024 604472
rect 399076 604460 399082 604512
rect 400858 604460 400864 604512
rect 400916 604500 400922 604512
rect 427354 604500 427360 604512
rect 400916 604472 427360 604500
rect 400916 604460 400922 604472
rect 427354 604460 427360 604472
rect 427412 604460 427418 604512
rect 428458 604460 428464 604512
rect 428516 604500 428522 604512
rect 455322 604500 455328 604512
rect 428516 604472 455328 604500
rect 428516 604460 428522 604472
rect 455322 604460 455328 604472
rect 455380 604460 455386 604512
rect 456150 604460 456156 604512
rect 456208 604500 456214 604512
rect 483014 604500 483020 604512
rect 456208 604472 483020 604500
rect 456208 604460 456214 604472
rect 483014 604460 483020 604472
rect 483072 604460 483078 604512
rect 485038 604460 485044 604512
rect 485096 604500 485102 604512
rect 511350 604500 511356 604512
rect 485096 604472 511356 604500
rect 485096 604460 485102 604472
rect 511350 604460 511356 604472
rect 511408 604460 511414 604512
rect 512638 604460 512644 604512
rect 512696 604500 512702 604512
rect 539318 604500 539324 604512
rect 512696 604472 539324 604500
rect 512696 604460 512702 604472
rect 539318 604460 539324 604472
rect 539376 604460 539382 604512
rect 540238 604460 540244 604512
rect 540296 604500 540302 604512
rect 567194 604500 567200 604512
rect 540296 604472 567200 604500
rect 540296 604460 540302 604472
rect 567194 604460 567200 604472
rect 567252 604460 567258 604512
rect 37918 602352 37924 602404
rect 37976 602392 37982 602404
rect 545758 602392 545764 602404
rect 37976 602364 545764 602392
rect 37976 602352 37982 602364
rect 545758 602352 545764 602364
rect 545816 602352 545822 602404
rect 35618 601672 35624 601724
rect 35676 601712 35682 601724
rect 36814 601712 36820 601724
rect 35676 601684 36820 601712
rect 35676 601672 35682 601684
rect 36814 601672 36820 601684
rect 36872 601672 36878 601724
rect 259730 584740 259736 584792
rect 259788 584780 259794 584792
rect 260190 584780 260196 584792
rect 259788 584752 260196 584780
rect 259788 584740 259794 584752
rect 260190 584740 260196 584752
rect 260248 584740 260254 584792
rect 148502 584400 148508 584452
rect 148560 584440 148566 584452
rect 155862 584440 155868 584452
rect 148560 584412 155868 584440
rect 148560 584400 148566 584412
rect 155862 584400 155868 584412
rect 155920 584400 155926 584452
rect 232682 584400 232688 584452
rect 232740 584440 232746 584452
rect 239766 584440 239772 584452
rect 232740 584412 239772 584440
rect 232740 584400 232746 584412
rect 239766 584400 239772 584412
rect 239824 584400 239830 584452
rect 428642 584400 428648 584452
rect 428700 584440 428706 584452
rect 435726 584440 435732 584452
rect 428700 584412 435732 584440
rect 428700 584400 428706 584412
rect 435726 584400 435732 584412
rect 435784 584400 435790 584452
rect 316770 584264 316776 584316
rect 316828 584304 316834 584316
rect 323854 584304 323860 584316
rect 316828 584276 323860 584304
rect 316828 584264 316834 584276
rect 323854 584264 323860 584276
rect 323912 584264 323918 584316
rect 512730 584264 512736 584316
rect 512788 584304 512794 584316
rect 519630 584304 519636 584316
rect 512788 584276 519636 584304
rect 512788 584264 512794 584276
rect 519630 584264 519636 584276
rect 519688 584264 519694 584316
rect 287698 584128 287704 584180
rect 287756 584168 287762 584180
rect 295702 584168 295708 584180
rect 287756 584140 295708 584168
rect 287756 584128 287762 584140
rect 295702 584128 295708 584140
rect 295760 584128 295766 584180
rect 483658 584128 483664 584180
rect 483716 584168 483722 584180
rect 491662 584168 491668 584180
rect 483716 584140 491668 584168
rect 483716 584128 483722 584140
rect 491662 584128 491668 584140
rect 491720 584128 491726 584180
rect 13722 583652 13728 583704
rect 13780 583692 13786 583704
rect 13780 583664 59952 583692
rect 13780 583652 13786 583664
rect 35618 583584 35624 583636
rect 35676 583624 35682 583636
rect 36998 583624 37004 583636
rect 35676 583596 37004 583624
rect 35676 583584 35682 583596
rect 36998 583584 37004 583596
rect 37056 583584 37062 583636
rect 42702 583584 42708 583636
rect 42760 583624 42766 583636
rect 42760 583596 45554 583624
rect 42760 583584 42766 583596
rect 45526 583488 45554 583596
rect 59924 583556 59952 583664
rect 63586 583652 63592 583704
rect 63644 583692 63650 583704
rect 64322 583692 64328 583704
rect 63644 583664 64328 583692
rect 63644 583652 63650 583664
rect 64322 583652 64328 583664
rect 64380 583652 64386 583704
rect 70302 583652 70308 583704
rect 70360 583692 70366 583704
rect 121454 583692 121460 583704
rect 70360 583664 121460 583692
rect 70360 583652 70366 583664
rect 121454 583652 121460 583664
rect 121512 583652 121518 583704
rect 126882 583652 126888 583704
rect 126940 583692 126946 583704
rect 178034 583692 178040 583704
rect 126940 583664 178040 583692
rect 126940 583652 126946 583664
rect 178034 583652 178040 583664
rect 178092 583652 178098 583704
rect 209682 583652 209688 583704
rect 209740 583692 209746 583704
rect 262214 583692 262220 583704
rect 209740 583664 262220 583692
rect 209740 583652 209746 583664
rect 262214 583652 262220 583664
rect 262272 583652 262278 583704
rect 266262 583652 266268 583704
rect 266320 583692 266326 583704
rect 317414 583692 317420 583704
rect 266320 583664 317420 583692
rect 266320 583652 266326 583664
rect 317414 583652 317420 583664
rect 317472 583652 317478 583704
rect 322842 583652 322848 583704
rect 322900 583692 322906 583704
rect 373994 583692 374000 583704
rect 322900 583664 374000 583692
rect 322900 583652 322906 583664
rect 373994 583652 374000 583664
rect 374052 583652 374058 583704
rect 405642 583652 405648 583704
rect 405700 583692 405706 583704
rect 458174 583692 458180 583704
rect 405700 583664 458180 583692
rect 405700 583652 405706 583664
rect 458174 583652 458180 583664
rect 458232 583652 458238 583704
rect 489822 583652 489828 583704
rect 489880 583692 489886 583704
rect 542354 583692 542360 583704
rect 489880 583664 542360 583692
rect 489880 583652 489886 583664
rect 542354 583652 542360 583664
rect 542412 583652 542418 583704
rect 93854 583624 93860 583636
rect 74506 583596 93860 583624
rect 66254 583556 66260 583568
rect 59924 583528 66260 583556
rect 66254 583516 66260 583528
rect 66312 583516 66318 583568
rect 74506 583488 74534 583596
rect 93854 583584 93860 583596
rect 93912 583584 93918 583636
rect 97902 583584 97908 583636
rect 97960 583624 97966 583636
rect 149054 583624 149060 583636
rect 97960 583596 149060 583624
rect 97960 583584 97966 583596
rect 149054 583584 149060 583596
rect 149112 583584 149118 583636
rect 154482 583584 154488 583636
rect 154540 583624 154546 583636
rect 205634 583624 205640 583636
rect 154540 583596 205640 583624
rect 154540 583584 154546 583596
rect 205634 583584 205640 583596
rect 205692 583584 205698 583636
rect 238662 583584 238668 583636
rect 238720 583624 238726 583636
rect 289814 583624 289820 583636
rect 238720 583596 289820 583624
rect 238720 583584 238726 583596
rect 289814 583584 289820 583596
rect 289872 583584 289878 583636
rect 293862 583584 293868 583636
rect 293920 583624 293926 583636
rect 293920 583596 335354 583624
rect 293920 583584 293926 583596
rect 182082 583516 182088 583568
rect 182140 583556 182146 583568
rect 233234 583556 233240 583568
rect 182140 583528 233240 583556
rect 182140 583516 182146 583528
rect 233234 583516 233240 583528
rect 233292 583516 233298 583568
rect 335326 583556 335354 583596
rect 343634 583584 343640 583636
rect 343692 583624 343698 583636
rect 345658 583624 345664 583636
rect 343692 583596 345664 583624
rect 343692 583584 343698 583596
rect 345658 583584 345664 583596
rect 345716 583584 345722 583636
rect 350442 583584 350448 583636
rect 350500 583624 350506 583636
rect 401594 583624 401600 583636
rect 350500 583596 401600 583624
rect 350500 583584 350506 583596
rect 401594 583584 401600 583596
rect 401652 583584 401658 583636
rect 427722 583584 427728 583636
rect 427780 583624 427786 583636
rect 428550 583624 428556 583636
rect 427780 583596 428556 583624
rect 427780 583584 427786 583596
rect 428550 583584 428556 583596
rect 428608 583584 428614 583636
rect 434622 583584 434628 583636
rect 434680 583624 434686 583636
rect 485774 583624 485780 583636
rect 434680 583596 485780 583624
rect 434680 583584 434686 583596
rect 485774 583584 485780 583596
rect 485832 583584 485838 583636
rect 518802 583584 518808 583636
rect 518860 583624 518866 583636
rect 569954 583624 569960 583636
rect 518860 583596 569960 583624
rect 518860 583584 518866 583596
rect 569954 583584 569960 583596
rect 570012 583584 570018 583636
rect 345014 583556 345020 583568
rect 335326 583528 345020 583556
rect 345014 583516 345020 583528
rect 345072 583516 345078 583568
rect 378042 583516 378048 583568
rect 378100 583556 378106 583568
rect 429194 583556 429200 583568
rect 378100 583528 429200 583556
rect 378100 583516 378106 583528
rect 429194 583516 429200 583528
rect 429252 583516 429258 583568
rect 462222 583516 462228 583568
rect 462280 583556 462286 583568
rect 513374 583556 513380 583568
rect 462280 583528 513380 583556
rect 462280 583516 462286 583528
rect 513374 583516 513380 583528
rect 513432 583516 513438 583568
rect 539502 583516 539508 583568
rect 539560 583556 539566 583568
rect 542998 583556 543004 583568
rect 539560 583528 543004 583556
rect 539560 583516 539566 583528
rect 542998 583516 543004 583528
rect 543056 583516 543062 583568
rect 45526 583460 74534 583488
rect 178678 580932 178684 580984
rect 178736 580972 178742 580984
rect 184014 580972 184020 580984
rect 178736 580944 184020 580972
rect 178736 580932 178742 580944
rect 184014 580932 184020 580944
rect 184072 580932 184078 580984
rect 374638 580932 374644 580984
rect 374696 580972 374702 580984
rect 379698 580972 379704 580984
rect 374696 580944 379704 580972
rect 374696 580932 374702 580944
rect 379698 580932 379704 580944
rect 379756 580932 379762 580984
rect 15194 580864 15200 580916
rect 15252 580904 15258 580916
rect 43990 580904 43996 580916
rect 15252 580876 43996 580904
rect 15252 580864 15258 580876
rect 43990 580864 43996 580876
rect 44048 580864 44054 580916
rect 71038 580864 71044 580916
rect 71096 580904 71102 580916
rect 567194 580904 567200 580916
rect 71096 580876 567200 580904
rect 71096 580864 71102 580876
rect 567194 580864 567200 580876
rect 567252 580864 567258 580916
rect 25682 580796 25688 580848
rect 25740 580836 25746 580848
rect 36906 580836 36912 580848
rect 25740 580808 36912 580836
rect 25740 580796 25746 580808
rect 36906 580796 36912 580808
rect 36964 580796 36970 580848
rect 53650 580796 53656 580848
rect 53708 580836 53714 580848
rect 66898 580836 66904 580848
rect 53708 580808 66904 580836
rect 53708 580796 53714 580808
rect 66898 580796 66904 580808
rect 66956 580796 66962 580848
rect 71866 580796 71872 580848
rect 71924 580836 71930 580848
rect 100018 580836 100024 580848
rect 71924 580808 100024 580836
rect 71924 580796 71930 580808
rect 100018 580796 100024 580808
rect 100076 580796 100082 580848
rect 127986 580836 127992 580848
rect 103486 580808 127992 580836
rect 42886 580728 42892 580780
rect 42944 580768 42950 580780
rect 72050 580768 72056 580780
rect 42944 580740 72056 580768
rect 42944 580728 42950 580740
rect 72050 580728 72056 580740
rect 72108 580728 72114 580780
rect 81986 580728 81992 580780
rect 82044 580768 82050 580780
rect 94498 580768 94504 580780
rect 82044 580740 94504 580768
rect 82044 580728 82050 580740
rect 94498 580728 94504 580740
rect 94556 580728 94562 580780
rect 99466 580728 99472 580780
rect 99524 580768 99530 580780
rect 103486 580768 103514 580808
rect 127986 580796 127992 580808
rect 128044 580796 128050 580848
rect 137646 580796 137652 580848
rect 137704 580836 137710 580848
rect 148410 580836 148416 580848
rect 137704 580808 148416 580836
rect 137704 580796 137710 580808
rect 148410 580796 148416 580808
rect 148468 580796 148474 580848
rect 165982 580796 165988 580848
rect 166040 580836 166046 580848
rect 177298 580836 177304 580848
rect 166040 580808 177304 580836
rect 166040 580796 166046 580808
rect 177298 580796 177304 580808
rect 177356 580796 177362 580848
rect 183646 580796 183652 580848
rect 183704 580836 183710 580848
rect 211706 580836 211712 580848
rect 183704 580808 211712 580836
rect 183704 580796 183710 580808
rect 211706 580796 211712 580808
rect 211764 580796 211770 580848
rect 222010 580796 222016 580848
rect 222068 580836 222074 580848
rect 232590 580836 232596 580848
rect 222068 580808 232596 580836
rect 222068 580796 222074 580808
rect 232590 580796 232596 580808
rect 232648 580796 232654 580848
rect 238846 580796 238852 580848
rect 238904 580836 238910 580848
rect 268010 580836 268016 580848
rect 238904 580808 268016 580836
rect 238904 580796 238910 580808
rect 268010 580796 268016 580808
rect 268068 580796 268074 580848
rect 277670 580796 277676 580848
rect 277728 580836 277734 580848
rect 289078 580836 289084 580848
rect 277728 580808 289084 580836
rect 277728 580796 277734 580808
rect 289078 580796 289084 580808
rect 289136 580796 289142 580848
rect 306006 580796 306012 580848
rect 306064 580836 306070 580848
rect 316678 580836 316684 580848
rect 306064 580808 316684 580836
rect 306064 580796 306070 580808
rect 316678 580796 316684 580808
rect 316736 580796 316742 580848
rect 323026 580796 323032 580848
rect 323084 580836 323090 580848
rect 352006 580836 352012 580848
rect 323084 580808 352012 580836
rect 323084 580796 323090 580808
rect 352006 580796 352012 580808
rect 352064 580796 352070 580848
rect 361666 580796 361672 580848
rect 361724 580836 361730 580848
rect 373258 580836 373264 580848
rect 361724 580808 373264 580836
rect 361724 580796 361730 580808
rect 373258 580796 373264 580808
rect 373316 580796 373322 580848
rect 379606 580796 379612 580848
rect 379664 580836 379670 580848
rect 408034 580836 408040 580848
rect 379664 580808 408040 580836
rect 379664 580796 379670 580808
rect 408034 580796 408040 580808
rect 408092 580796 408098 580848
rect 417694 580796 417700 580848
rect 417752 580836 417758 580848
rect 428458 580836 428464 580848
rect 417752 580808 428464 580836
rect 417752 580796 417758 580808
rect 428458 580796 428464 580808
rect 428516 580796 428522 580848
rect 434806 580796 434812 580848
rect 434864 580836 434870 580848
rect 463694 580836 463700 580848
rect 434864 580808 463700 580836
rect 434864 580796 434870 580808
rect 463694 580796 463700 580808
rect 463752 580796 463758 580848
rect 473998 580796 474004 580848
rect 474056 580836 474062 580848
rect 485038 580836 485044 580848
rect 474056 580808 485044 580836
rect 474056 580796 474062 580808
rect 485038 580796 485044 580808
rect 485096 580796 485102 580848
rect 501690 580796 501696 580848
rect 501748 580836 501754 580848
rect 512638 580836 512644 580848
rect 501748 580808 512644 580836
rect 501748 580796 501754 580808
rect 512638 580796 512644 580808
rect 512696 580796 512702 580848
rect 518986 580796 518992 580848
rect 519044 580836 519050 580848
rect 547874 580836 547880 580848
rect 519044 580808 547880 580836
rect 519044 580796 519050 580808
rect 547874 580796 547880 580808
rect 547932 580796 547938 580848
rect 99524 580740 103514 580768
rect 99524 580728 99530 580740
rect 109678 580728 109684 580780
rect 109736 580768 109742 580780
rect 120718 580768 120724 580780
rect 109736 580740 120724 580768
rect 109736 580728 109742 580740
rect 120718 580728 120724 580740
rect 120776 580728 120782 580780
rect 193674 580728 193680 580780
rect 193732 580768 193738 580780
rect 204898 580768 204904 580780
rect 193732 580740 204904 580768
rect 193732 580728 193738 580740
rect 204898 580728 204904 580740
rect 204956 580728 204962 580780
rect 249702 580728 249708 580780
rect 249760 580768 249766 580780
rect 260098 580768 260104 580780
rect 249760 580740 260104 580768
rect 249760 580728 249766 580740
rect 260098 580728 260104 580740
rect 260156 580728 260162 580780
rect 333698 580728 333704 580780
rect 333756 580768 333762 580780
rect 344278 580768 344284 580780
rect 333756 580740 344284 580768
rect 333756 580728 333762 580740
rect 344278 580728 344284 580740
rect 344336 580728 344342 580780
rect 390002 580728 390008 580780
rect 390060 580768 390066 580780
rect 400858 580768 400864 580780
rect 390060 580740 400864 580768
rect 390060 580728 390066 580740
rect 400858 580728 400864 580740
rect 400916 580728 400922 580780
rect 445662 580728 445668 580780
rect 445720 580768 445726 580780
rect 456150 580768 456156 580780
rect 445720 580740 456156 580768
rect 445720 580728 445726 580740
rect 456150 580728 456156 580740
rect 456208 580728 456214 580780
rect 529658 580728 529664 580780
rect 529716 580768 529722 580780
rect 540238 580768 540244 580780
rect 529716 580740 540244 580768
rect 529716 580728 529722 580740
rect 540238 580728 540244 580740
rect 540296 580728 540302 580780
rect 36722 580660 36728 580712
rect 36780 580700 36786 580712
rect 557534 580700 557540 580712
rect 36780 580672 557540 580700
rect 36780 580660 36786 580672
rect 557534 580660 557540 580672
rect 557592 580660 557598 580712
rect 3234 579708 3240 579760
rect 3292 579748 3298 579760
rect 7558 579748 7564 579760
rect 3292 579720 7564 579748
rect 3292 579708 3298 579720
rect 7558 579708 7564 579720
rect 7616 579708 7622 579760
rect 16022 578892 16028 578944
rect 16080 578932 16086 578944
rect 547874 578932 547880 578944
rect 16080 578904 547880 578932
rect 16080 578892 16086 578904
rect 547874 578892 547880 578904
rect 547932 578892 547938 578944
rect 25682 578416 25688 578468
rect 25740 578456 25746 578468
rect 71038 578456 71044 578468
rect 25740 578428 71044 578456
rect 25740 578416 25746 578428
rect 71038 578416 71044 578428
rect 71096 578416 71102 578468
rect 296346 578416 296352 578468
rect 296404 578456 296410 578468
rect 316770 578456 316776 578468
rect 296404 578428 316776 578456
rect 296404 578416 296410 578428
rect 316770 578416 316776 578428
rect 316828 578416 316834 578468
rect 408034 578416 408040 578468
rect 408092 578456 408098 578468
rect 428642 578456 428648 578468
rect 408092 578428 428648 578456
rect 408092 578416 408098 578428
rect 428642 578416 428648 578428
rect 428700 578416 428706 578468
rect 492030 578416 492036 578468
rect 492088 578456 492094 578468
rect 512730 578456 512736 578468
rect 492088 578428 512736 578456
rect 492088 578416 492094 578428
rect 512730 578416 512736 578428
rect 512788 578416 512794 578468
rect 36906 578348 36912 578400
rect 36964 578388 36970 578400
rect 53650 578388 53656 578400
rect 36964 578360 53656 578388
rect 36964 578348 36970 578360
rect 53650 578348 53656 578360
rect 53708 578348 53714 578400
rect 148410 578348 148416 578400
rect 148468 578388 148474 578400
rect 165614 578388 165620 578400
rect 148468 578360 165620 578388
rect 148468 578348 148474 578360
rect 165614 578348 165620 578360
rect 165672 578348 165678 578400
rect 175458 578348 175464 578400
rect 175516 578388 175522 578400
rect 193674 578388 193680 578400
rect 175516 578360 193680 578388
rect 175516 578348 175522 578360
rect 193674 578348 193680 578360
rect 193732 578348 193738 578400
rect 203518 578348 203524 578400
rect 203576 578388 203582 578400
rect 221366 578388 221372 578400
rect 203576 578360 221372 578388
rect 203576 578348 203582 578360
rect 221366 578348 221372 578360
rect 221424 578348 221430 578400
rect 232498 578348 232504 578400
rect 232556 578388 232562 578400
rect 249702 578388 249708 578400
rect 232556 578360 249708 578388
rect 232556 578348 232562 578360
rect 249702 578348 249708 578360
rect 249760 578348 249766 578400
rect 260190 578348 260196 578400
rect 260248 578388 260254 578400
rect 277670 578388 277676 578400
rect 260248 578360 277676 578388
rect 260248 578348 260254 578360
rect 277670 578348 277676 578360
rect 277728 578348 277734 578400
rect 287514 578348 287520 578400
rect 287572 578388 287578 578400
rect 305362 578388 305368 578400
rect 287572 578360 305368 578388
rect 287572 578348 287578 578360
rect 305362 578348 305368 578360
rect 305420 578348 305426 578400
rect 345658 578348 345664 578400
rect 345716 578388 345722 578400
rect 361666 578388 361672 578400
rect 345716 578360 361672 578388
rect 345716 578348 345722 578360
rect 361666 578348 361672 578360
rect 361724 578348 361730 578400
rect 371510 578348 371516 578400
rect 371568 578388 371574 578400
rect 389358 578388 389364 578400
rect 371568 578360 389364 578388
rect 371568 578348 371574 578360
rect 389358 578348 389364 578360
rect 389416 578348 389422 578400
rect 399478 578348 399484 578400
rect 399536 578388 399542 578400
rect 417694 578388 417700 578400
rect 399536 578360 417700 578388
rect 399536 578348 399542 578360
rect 417694 578348 417700 578360
rect 417752 578348 417758 578400
rect 456150 578348 456156 578400
rect 456208 578388 456214 578400
rect 473538 578388 473544 578400
rect 456208 578360 473544 578388
rect 456208 578348 456214 578360
rect 473538 578348 473544 578360
rect 473596 578348 473602 578400
rect 483474 578348 483480 578400
rect 483532 578388 483538 578400
rect 501690 578388 501696 578400
rect 483532 578360 501696 578388
rect 483532 578348 483538 578360
rect 501690 578348 501696 578360
rect 501748 578348 501754 578400
rect 36998 578280 37004 578332
rect 37056 578320 37062 578332
rect 63310 578320 63316 578332
rect 37056 578292 63316 578320
rect 37056 578280 37062 578292
rect 63310 578280 63316 578292
rect 63368 578280 63374 578332
rect 64322 578280 64328 578332
rect 64380 578320 64386 578332
rect 81434 578320 81440 578332
rect 64380 578292 81440 578320
rect 64380 578280 64386 578292
rect 81434 578280 81440 578292
rect 81492 578280 81498 578332
rect 91462 578280 91468 578332
rect 91520 578320 91526 578332
rect 109678 578320 109684 578332
rect 91520 578292 109684 578320
rect 91520 578280 91526 578292
rect 109678 578280 109684 578292
rect 109736 578280 109742 578332
rect 119430 578280 119436 578332
rect 119488 578320 119494 578332
rect 137646 578320 137652 578332
rect 119488 578292 137652 578320
rect 119488 578280 119494 578292
rect 137646 578280 137652 578292
rect 137704 578280 137710 578332
rect 156322 578280 156328 578332
rect 156380 578320 156386 578332
rect 178678 578320 178684 578332
rect 156380 578292 178684 578320
rect 156380 578280 156386 578292
rect 178678 578280 178684 578292
rect 178736 578280 178742 578332
rect 212258 578280 212264 578332
rect 212316 578320 212322 578332
rect 232682 578320 232688 578332
rect 212316 578292 232688 578320
rect 212316 578280 212322 578292
rect 232682 578280 232688 578292
rect 232740 578280 232746 578332
rect 268010 578280 268016 578332
rect 268068 578320 268074 578332
rect 287698 578320 287704 578332
rect 268068 578292 287704 578320
rect 268068 578280 268074 578292
rect 287698 578280 287704 578292
rect 287756 578280 287762 578332
rect 315482 578280 315488 578332
rect 315540 578320 315546 578332
rect 333698 578320 333704 578332
rect 315540 578292 333704 578320
rect 315540 578280 315546 578292
rect 333698 578280 333704 578292
rect 333756 578280 333762 578332
rect 352006 578280 352012 578332
rect 352064 578320 352070 578332
rect 374638 578320 374644 578332
rect 352064 578292 374644 578320
rect 352064 578280 352070 578292
rect 374638 578280 374644 578292
rect 374696 578280 374702 578332
rect 428458 578280 428464 578332
rect 428516 578320 428522 578332
rect 445662 578320 445668 578332
rect 428516 578292 445668 578320
rect 428516 578280 428522 578292
rect 445662 578280 445668 578292
rect 445720 578280 445726 578332
rect 464338 578280 464344 578332
rect 464396 578320 464402 578332
rect 483658 578320 483664 578332
rect 464396 578292 483664 578320
rect 464396 578280 464402 578292
rect 483658 578280 483664 578292
rect 483716 578280 483722 578332
rect 511442 578280 511448 578332
rect 511500 578320 511506 578332
rect 529658 578320 529664 578332
rect 511500 578292 529664 578320
rect 511500 578280 511506 578292
rect 529658 578280 529664 578292
rect 529716 578280 529722 578332
rect 542998 578280 543004 578332
rect 543056 578320 543062 578332
rect 557534 578320 557540 578332
rect 543056 578292 557540 578320
rect 543056 578280 543062 578292
rect 557534 578280 557540 578292
rect 557592 578280 557598 578332
rect 69658 578212 69664 578264
rect 69716 578252 69722 578264
rect 91094 578252 91100 578264
rect 69716 578224 91100 578252
rect 69716 578212 69722 578224
rect 91094 578212 91100 578224
rect 91152 578212 91158 578264
rect 94498 578212 94504 578264
rect 94556 578252 94562 578264
rect 119338 578252 119344 578264
rect 94556 578224 119344 578252
rect 94556 578212 94562 578224
rect 119338 578212 119344 578224
rect 119396 578212 119402 578264
rect 120718 578212 120724 578264
rect 120776 578252 120782 578264
rect 147306 578252 147312 578264
rect 120776 578224 147312 578252
rect 120776 578212 120782 578224
rect 147306 578212 147312 578224
rect 147364 578212 147370 578264
rect 148318 578212 148324 578264
rect 148376 578252 148382 578264
rect 175274 578252 175280 578264
rect 148376 578224 175280 578252
rect 148376 578212 148382 578224
rect 175274 578212 175280 578224
rect 175332 578212 175338 578264
rect 177298 578212 177304 578264
rect 177356 578252 177362 578264
rect 203334 578252 203340 578264
rect 177356 578224 203340 578252
rect 177356 578212 177362 578224
rect 203334 578212 203340 578224
rect 203392 578212 203398 578264
rect 204898 578212 204904 578264
rect 204956 578252 204962 578264
rect 231026 578252 231032 578264
rect 204956 578224 231032 578252
rect 204956 578212 204962 578224
rect 231026 578212 231032 578224
rect 231084 578212 231090 578264
rect 232590 578212 232596 578264
rect 232648 578252 232654 578264
rect 259362 578252 259368 578264
rect 232648 578224 259368 578252
rect 232648 578212 232654 578224
rect 259362 578212 259368 578224
rect 259420 578212 259426 578264
rect 260098 578212 260104 578264
rect 260156 578252 260162 578264
rect 287330 578252 287336 578264
rect 260156 578224 287336 578252
rect 260156 578212 260162 578224
rect 287330 578212 287336 578224
rect 287388 578212 287394 578264
rect 289078 578212 289084 578264
rect 289136 578252 289142 578264
rect 315022 578252 315028 578264
rect 289136 578224 315028 578252
rect 289136 578212 289142 578224
rect 315022 578212 315028 578224
rect 315080 578212 315086 578264
rect 316678 578212 316684 578264
rect 316736 578252 316742 578264
rect 343358 578252 343364 578264
rect 316736 578224 343364 578252
rect 316736 578212 316742 578224
rect 343358 578212 343364 578224
rect 343416 578212 343422 578264
rect 344278 578212 344284 578264
rect 344336 578252 344342 578264
rect 371326 578252 371332 578264
rect 344336 578224 371332 578252
rect 344336 578212 344342 578224
rect 371326 578212 371332 578224
rect 371384 578212 371390 578264
rect 373258 578212 373264 578264
rect 373316 578252 373322 578264
rect 399018 578252 399024 578264
rect 373316 578224 399024 578252
rect 373316 578212 373322 578224
rect 399018 578212 399024 578224
rect 399076 578212 399082 578264
rect 400858 578212 400864 578264
rect 400916 578252 400922 578264
rect 427354 578252 427360 578264
rect 400916 578224 427360 578252
rect 400916 578212 400922 578224
rect 427354 578212 427360 578224
rect 427412 578212 427418 578264
rect 428550 578212 428556 578264
rect 428608 578252 428614 578264
rect 455322 578252 455328 578264
rect 428608 578224 455328 578252
rect 428608 578212 428614 578224
rect 455322 578212 455328 578224
rect 455380 578212 455386 578264
rect 456058 578212 456064 578264
rect 456116 578252 456122 578264
rect 483198 578252 483204 578264
rect 456116 578224 483204 578252
rect 456116 578212 456122 578224
rect 483198 578212 483204 578224
rect 483256 578212 483262 578264
rect 485038 578212 485044 578264
rect 485096 578252 485102 578264
rect 511350 578252 511356 578264
rect 485096 578224 511356 578252
rect 485096 578212 485102 578224
rect 511350 578212 511356 578224
rect 511408 578212 511414 578264
rect 512638 578212 512644 578264
rect 512696 578252 512702 578264
rect 539318 578252 539324 578264
rect 512696 578224 539324 578252
rect 512696 578212 512702 578224
rect 539318 578212 539324 578224
rect 539376 578212 539382 578264
rect 540238 578212 540244 578264
rect 540296 578252 540302 578264
rect 567194 578252 567200 578264
rect 540296 578224 567200 578252
rect 540296 578212 540302 578224
rect 567194 578212 567200 578224
rect 567252 578212 567258 578264
rect 37918 576104 37924 576156
rect 37976 576144 37982 576156
rect 545758 576144 545764 576156
rect 37976 576116 545764 576144
rect 37976 576104 37982 576116
rect 545758 576104 545764 576116
rect 545816 576104 545822 576156
rect 35618 575424 35624 575476
rect 35676 575464 35682 575476
rect 36722 575464 36728 575476
rect 35676 575436 36728 575464
rect 35676 575424 35682 575436
rect 36722 575424 36728 575436
rect 36780 575424 36786 575476
rect 147674 562300 147680 562352
rect 147732 562340 147738 562352
rect 148410 562340 148416 562352
rect 147732 562312 148416 562340
rect 147732 562300 147738 562312
rect 148410 562300 148416 562312
rect 148468 562300 148474 562352
rect 259730 562300 259736 562352
rect 259788 562340 259794 562352
rect 260190 562340 260196 562352
rect 259788 562312 260196 562340
rect 259788 562300 259794 562312
rect 260190 562300 260196 562312
rect 260248 562300 260254 562352
rect 455690 562300 455696 562352
rect 455748 562340 455754 562352
rect 456150 562340 456156 562352
rect 455748 562312 456156 562340
rect 455748 562300 455754 562312
rect 456150 562300 456156 562312
rect 456208 562300 456214 562352
rect 287698 558832 287704 558884
rect 287756 558872 287762 558884
rect 295702 558872 295708 558884
rect 287756 558844 295708 558872
rect 287756 558832 287762 558844
rect 295702 558832 295708 558844
rect 295760 558832 295766 558884
rect 316770 558832 316776 558884
rect 316828 558872 316834 558884
rect 323670 558872 323676 558884
rect 316828 558844 323676 558872
rect 316828 558832 316834 558844
rect 323670 558832 323676 558844
rect 323728 558832 323734 558884
rect 63586 558288 63592 558340
rect 63644 558328 63650 558340
rect 64322 558328 64328 558340
rect 63644 558300 64328 558328
rect 63644 558288 63650 558300
rect 64322 558288 64328 558300
rect 64380 558288 64386 558340
rect 232682 558152 232688 558204
rect 232740 558192 232746 558204
rect 239766 558192 239772 558204
rect 232740 558164 239772 558192
rect 232740 558152 232746 558164
rect 239766 558152 239772 558164
rect 239824 558152 239830 558204
rect 428642 558152 428648 558204
rect 428700 558192 428706 558204
rect 435726 558192 435732 558204
rect 428700 558164 435732 558192
rect 428700 558152 428706 558164
rect 435726 558152 435732 558164
rect 435784 558152 435790 558204
rect 483658 558152 483664 558204
rect 483716 558192 483722 558204
rect 491662 558192 491668 558204
rect 483716 558164 491668 558192
rect 483716 558152 483722 558164
rect 491662 558152 491668 558164
rect 491720 558152 491726 558204
rect 512730 557608 512736 557660
rect 512788 557648 512794 557660
rect 519630 557648 519636 557660
rect 512788 557620 519636 557648
rect 512788 557608 512794 557620
rect 519630 557608 519636 557620
rect 519688 557608 519694 557660
rect 13722 557472 13728 557524
rect 13780 557512 13786 557524
rect 66254 557512 66260 557524
rect 13780 557484 66260 557512
rect 13780 557472 13786 557484
rect 66254 557472 66260 557484
rect 66312 557472 66318 557524
rect 97902 557472 97908 557524
rect 97960 557512 97966 557524
rect 149054 557512 149060 557524
rect 97960 557484 149060 557512
rect 97960 557472 97966 557484
rect 149054 557472 149060 557484
rect 149112 557472 149118 557524
rect 154482 557472 154488 557524
rect 154540 557512 154546 557524
rect 205634 557512 205640 557524
rect 154540 557484 205640 557512
rect 154540 557472 154546 557484
rect 205634 557472 205640 557484
rect 205692 557472 205698 557524
rect 209682 557472 209688 557524
rect 209740 557512 209746 557524
rect 262214 557512 262220 557524
rect 209740 557484 262220 557512
rect 209740 557472 209746 557484
rect 262214 557472 262220 557484
rect 262272 557472 262278 557524
rect 266262 557472 266268 557524
rect 266320 557512 266326 557524
rect 317414 557512 317420 557524
rect 266320 557484 317420 557512
rect 266320 557472 266326 557484
rect 317414 557472 317420 557484
rect 317472 557472 317478 557524
rect 322842 557472 322848 557524
rect 322900 557512 322906 557524
rect 373994 557512 374000 557524
rect 322900 557484 374000 557512
rect 322900 557472 322906 557484
rect 373994 557472 374000 557484
rect 374052 557472 374058 557524
rect 405642 557472 405648 557524
rect 405700 557512 405706 557524
rect 458174 557512 458180 557524
rect 405700 557484 458180 557512
rect 405700 557472 405706 557484
rect 458174 557472 458180 557484
rect 458232 557472 458238 557524
rect 489822 557472 489828 557524
rect 489880 557512 489886 557524
rect 542354 557512 542360 557524
rect 489880 557484 542360 557512
rect 489880 557472 489886 557484
rect 542354 557472 542360 557484
rect 542412 557472 542418 557524
rect 35618 557404 35624 557456
rect 35676 557444 35682 557456
rect 36906 557444 36912 557456
rect 35676 557416 36912 557444
rect 35676 557404 35682 557416
rect 36906 557404 36912 557416
rect 36964 557404 36970 557456
rect 42702 557404 42708 557456
rect 42760 557444 42766 557456
rect 93854 557444 93860 557456
rect 42760 557416 93860 557444
rect 42760 557404 42766 557416
rect 93854 557404 93860 557416
rect 93912 557404 93918 557456
rect 126882 557404 126888 557456
rect 126940 557444 126946 557456
rect 178034 557444 178040 557456
rect 126940 557416 178040 557444
rect 126940 557404 126946 557416
rect 178034 557404 178040 557416
rect 178092 557404 178098 557456
rect 182082 557404 182088 557456
rect 182140 557444 182146 557456
rect 233234 557444 233240 557456
rect 182140 557416 233240 557444
rect 182140 557404 182146 557416
rect 233234 557404 233240 557416
rect 233292 557404 233298 557456
rect 238662 557404 238668 557456
rect 238720 557444 238726 557456
rect 289814 557444 289820 557456
rect 238720 557416 289820 557444
rect 238720 557404 238726 557416
rect 289814 557404 289820 557416
rect 289872 557404 289878 557456
rect 293862 557404 293868 557456
rect 293920 557444 293926 557456
rect 293920 557416 335354 557444
rect 293920 557404 293926 557416
rect 70302 557336 70308 557388
rect 70360 557376 70366 557388
rect 121454 557376 121460 557388
rect 70360 557348 121460 557376
rect 70360 557336 70366 557348
rect 121454 557336 121460 557348
rect 121512 557336 121518 557388
rect 335326 557376 335354 557416
rect 343542 557404 343548 557456
rect 343600 557444 343606 557456
rect 345658 557444 345664 557456
rect 343600 557416 345664 557444
rect 343600 557404 343606 557416
rect 345658 557404 345664 557416
rect 345716 557404 345722 557456
rect 350442 557404 350448 557456
rect 350500 557444 350506 557456
rect 401594 557444 401600 557456
rect 350500 557416 401600 557444
rect 350500 557404 350506 557416
rect 401594 557404 401600 557416
rect 401652 557404 401658 557456
rect 434622 557404 434628 557456
rect 434680 557444 434686 557456
rect 485774 557444 485780 557456
rect 434680 557416 485780 557444
rect 434680 557404 434686 557416
rect 485774 557404 485780 557416
rect 485832 557404 485838 557456
rect 518802 557404 518808 557456
rect 518860 557444 518866 557456
rect 569954 557444 569960 557456
rect 518860 557416 569960 557444
rect 518860 557404 518866 557416
rect 569954 557404 569960 557416
rect 570012 557404 570018 557456
rect 345014 557376 345020 557388
rect 335326 557348 345020 557376
rect 345014 557336 345020 557348
rect 345072 557336 345078 557388
rect 378042 557336 378048 557388
rect 378100 557376 378106 557388
rect 429194 557376 429200 557388
rect 378100 557348 429200 557376
rect 378100 557336 378106 557348
rect 429194 557336 429200 557348
rect 429252 557336 429258 557388
rect 462222 557336 462228 557388
rect 462280 557376 462286 557388
rect 513374 557376 513380 557388
rect 462280 557348 513380 557376
rect 462280 557336 462286 557348
rect 513374 557336 513380 557348
rect 513432 557336 513438 557388
rect 42886 554684 42892 554736
rect 42944 554724 42950 554736
rect 72050 554724 72056 554736
rect 42944 554696 45554 554724
rect 42944 554684 42950 554696
rect 15194 554616 15200 554668
rect 15252 554656 15258 554668
rect 43990 554656 43996 554668
rect 15252 554628 43996 554656
rect 15252 554616 15258 554628
rect 43990 554616 43996 554628
rect 44048 554616 44054 554668
rect 45526 554656 45554 554696
rect 64846 554696 72056 554724
rect 64846 554656 64874 554696
rect 72050 554684 72056 554696
rect 72108 554684 72114 554736
rect 99466 554684 99472 554736
rect 99524 554724 99530 554736
rect 99524 554696 103514 554724
rect 99524 554684 99530 554696
rect 45526 554628 64874 554656
rect 71866 554616 71872 554668
rect 71924 554656 71930 554668
rect 100018 554656 100024 554668
rect 71924 554628 100024 554656
rect 71924 554616 71930 554628
rect 100018 554616 100024 554628
rect 100076 554616 100082 554668
rect 103486 554656 103514 554696
rect 127066 554684 127072 554736
rect 127124 554724 127130 554736
rect 127124 554696 132494 554724
rect 127124 554684 127130 554696
rect 127986 554656 127992 554668
rect 103486 554628 127992 554656
rect 127986 554616 127992 554628
rect 128044 554616 128050 554668
rect 132466 554656 132494 554696
rect 183646 554684 183652 554736
rect 183704 554724 183710 554736
rect 183704 554696 190454 554724
rect 183704 554684 183710 554696
rect 156046 554656 156052 554668
rect 132466 554628 156052 554656
rect 156046 554616 156052 554628
rect 156104 554616 156110 554668
rect 165982 554616 165988 554668
rect 166040 554656 166046 554668
rect 177298 554656 177304 554668
rect 166040 554628 177304 554656
rect 166040 554616 166046 554628
rect 177298 554616 177304 554628
rect 177356 554616 177362 554668
rect 178678 554616 178684 554668
rect 178736 554656 178742 554668
rect 184014 554656 184020 554668
rect 178736 554628 184020 554656
rect 178736 554616 178742 554628
rect 184014 554616 184020 554628
rect 184072 554616 184078 554668
rect 190426 554656 190454 554696
rect 374638 554684 374644 554736
rect 374696 554724 374702 554736
rect 379698 554724 379704 554736
rect 374696 554696 379704 554724
rect 374696 554684 374702 554696
rect 379698 554684 379704 554696
rect 379756 554684 379762 554736
rect 539318 554684 539324 554736
rect 539376 554724 539382 554736
rect 542998 554724 543004 554736
rect 539376 554696 543004 554724
rect 539376 554684 539382 554696
rect 542998 554684 543004 554696
rect 543056 554684 543062 554736
rect 211706 554656 211712 554668
rect 190426 554628 211712 554656
rect 211706 554616 211712 554628
rect 211764 554616 211770 554668
rect 222010 554616 222016 554668
rect 222068 554656 222074 554668
rect 232590 554656 232596 554668
rect 222068 554628 232596 554656
rect 222068 554616 222074 554628
rect 232590 554616 232596 554628
rect 232648 554616 232654 554668
rect 249702 554616 249708 554668
rect 249760 554656 249766 554668
rect 260098 554656 260104 554668
rect 249760 554628 260104 554656
rect 249760 554616 249766 554628
rect 260098 554616 260104 554628
rect 260156 554616 260162 554668
rect 261478 554616 261484 554668
rect 261536 554656 261542 554668
rect 567194 554656 567200 554668
rect 261536 554628 567200 554656
rect 261536 554616 261542 554628
rect 567194 554616 567200 554628
rect 567252 554616 567258 554668
rect 25682 554548 25688 554600
rect 25740 554588 25746 554600
rect 36998 554588 37004 554600
rect 25740 554560 37004 554588
rect 25740 554548 25746 554560
rect 36998 554548 37004 554560
rect 37056 554548 37062 554600
rect 53650 554548 53656 554600
rect 53708 554588 53714 554600
rect 69658 554588 69664 554600
rect 53708 554560 69664 554588
rect 53708 554548 53714 554560
rect 69658 554548 69664 554560
rect 69716 554548 69722 554600
rect 81986 554548 81992 554600
rect 82044 554588 82050 554600
rect 94498 554588 94504 554600
rect 82044 554560 94504 554588
rect 82044 554548 82050 554560
rect 94498 554548 94504 554560
rect 94556 554548 94562 554600
rect 109678 554548 109684 554600
rect 109736 554588 109742 554600
rect 120718 554588 120724 554600
rect 109736 554560 120724 554588
rect 109736 554548 109742 554560
rect 120718 554548 120724 554560
rect 120776 554548 120782 554600
rect 137646 554548 137652 554600
rect 137704 554588 137710 554600
rect 148318 554588 148324 554600
rect 137704 554560 148324 554588
rect 137704 554548 137710 554560
rect 148318 554548 148324 554560
rect 148376 554548 148382 554600
rect 193674 554548 193680 554600
rect 193732 554588 193738 554600
rect 204898 554588 204904 554600
rect 193732 554560 204904 554588
rect 193732 554548 193738 554560
rect 204898 554548 204904 554560
rect 204956 554548 204962 554600
rect 238846 554548 238852 554600
rect 238904 554588 238910 554600
rect 268010 554588 268016 554600
rect 238904 554560 268016 554588
rect 238904 554548 238910 554560
rect 268010 554548 268016 554560
rect 268068 554548 268074 554600
rect 277670 554548 277676 554600
rect 277728 554588 277734 554600
rect 289078 554588 289084 554600
rect 277728 554560 289084 554588
rect 277728 554548 277734 554560
rect 289078 554548 289084 554560
rect 289136 554548 289142 554600
rect 306006 554548 306012 554600
rect 306064 554588 306070 554600
rect 316678 554588 316684 554600
rect 306064 554560 316684 554588
rect 306064 554548 306070 554560
rect 316678 554548 316684 554560
rect 316736 554548 316742 554600
rect 323026 554548 323032 554600
rect 323084 554588 323090 554600
rect 352006 554588 352012 554600
rect 323084 554560 352012 554588
rect 323084 554548 323090 554560
rect 352006 554548 352012 554560
rect 352064 554548 352070 554600
rect 361666 554548 361672 554600
rect 361724 554588 361730 554600
rect 373258 554588 373264 554600
rect 361724 554560 373264 554588
rect 361724 554548 361730 554560
rect 373258 554548 373264 554560
rect 373316 554548 373322 554600
rect 379606 554548 379612 554600
rect 379664 554588 379670 554600
rect 408034 554588 408040 554600
rect 379664 554560 408040 554588
rect 379664 554548 379670 554560
rect 408034 554548 408040 554560
rect 408092 554548 408098 554600
rect 417694 554548 417700 554600
rect 417752 554588 417758 554600
rect 428550 554588 428556 554600
rect 417752 554560 428556 554588
rect 417752 554548 417758 554560
rect 428550 554548 428556 554560
rect 428608 554548 428614 554600
rect 434806 554548 434812 554600
rect 434864 554588 434870 554600
rect 463694 554588 463700 554600
rect 434864 554560 463700 554588
rect 434864 554548 434870 554560
rect 463694 554548 463700 554560
rect 463752 554548 463758 554600
rect 473998 554548 474004 554600
rect 474056 554588 474062 554600
rect 485038 554588 485044 554600
rect 474056 554560 485044 554588
rect 474056 554548 474062 554560
rect 485038 554548 485044 554560
rect 485096 554548 485102 554600
rect 501690 554548 501696 554600
rect 501748 554588 501754 554600
rect 512638 554588 512644 554600
rect 501748 554560 512644 554588
rect 501748 554548 501754 554560
rect 512638 554548 512644 554560
rect 512696 554548 512702 554600
rect 518986 554548 518992 554600
rect 519044 554588 519050 554600
rect 547874 554588 547880 554600
rect 519044 554560 547880 554588
rect 519044 554548 519050 554560
rect 547874 554548 547880 554560
rect 547932 554548 547938 554600
rect 333698 554480 333704 554532
rect 333756 554520 333762 554532
rect 344278 554520 344284 554532
rect 333756 554492 344284 554520
rect 333756 554480 333762 554492
rect 344278 554480 344284 554492
rect 344336 554480 344342 554532
rect 390002 554480 390008 554532
rect 390060 554520 390066 554532
rect 400858 554520 400864 554532
rect 390060 554492 400864 554520
rect 390060 554480 390066 554492
rect 400858 554480 400864 554492
rect 400916 554480 400922 554532
rect 445662 554480 445668 554532
rect 445720 554520 445726 554532
rect 456058 554520 456064 554532
rect 445720 554492 456064 554520
rect 445720 554480 445726 554492
rect 456058 554480 456064 554492
rect 456116 554480 456122 554532
rect 529658 554480 529664 554532
rect 529716 554520 529722 554532
rect 540238 554520 540244 554532
rect 529716 554492 540244 554520
rect 529716 554480 529722 554492
rect 540238 554480 540244 554492
rect 540296 554480 540302 554532
rect 36814 554412 36820 554464
rect 36872 554452 36878 554464
rect 557534 554452 557540 554464
rect 36872 554424 557540 554452
rect 36872 554412 36878 554424
rect 557534 554412 557540 554424
rect 557592 554412 557598 554464
rect 16022 551284 16028 551336
rect 16080 551324 16086 551336
rect 547874 551324 547880 551336
rect 16080 551296 547880 551324
rect 16080 551284 16086 551296
rect 547874 551284 547880 551296
rect 547932 551284 547938 551336
rect 25682 550876 25688 550928
rect 25740 550916 25746 550928
rect 261478 550916 261484 550928
rect 25740 550888 261484 550916
rect 25740 550876 25746 550888
rect 261478 550876 261484 550888
rect 261536 550876 261542 550928
rect 148318 550808 148324 550860
rect 148376 550848 148382 550860
rect 165706 550848 165712 550860
rect 148376 550820 165712 550848
rect 148376 550808 148382 550820
rect 165706 550808 165712 550820
rect 165764 550808 165770 550860
rect 175458 550808 175464 550860
rect 175516 550848 175522 550860
rect 193674 550848 193680 550860
rect 175516 550820 193680 550848
rect 175516 550808 175522 550820
rect 193674 550808 193680 550820
rect 193732 550808 193738 550860
rect 203518 550808 203524 550860
rect 203576 550848 203582 550860
rect 221366 550848 221372 550860
rect 203576 550820 221372 550848
rect 203576 550808 203582 550820
rect 221366 550808 221372 550820
rect 221424 550808 221430 550860
rect 296346 550808 296352 550860
rect 296404 550848 296410 550860
rect 316770 550848 316776 550860
rect 296404 550820 316776 550848
rect 296404 550808 296410 550820
rect 316770 550808 316776 550820
rect 316828 550808 316834 550860
rect 408034 550808 408040 550860
rect 408092 550848 408098 550860
rect 428642 550848 428648 550860
rect 408092 550820 428648 550848
rect 408092 550808 408098 550820
rect 428642 550808 428648 550820
rect 428700 550808 428706 550860
rect 492030 550808 492036 550860
rect 492088 550848 492094 550860
rect 512730 550848 512736 550860
rect 492088 550820 512736 550848
rect 492088 550808 492094 550820
rect 512730 550808 512736 550820
rect 512788 550808 512794 550860
rect 36814 550740 36820 550792
rect 36872 550780 36878 550792
rect 53650 550780 53656 550792
rect 36872 550752 53656 550780
rect 36872 550740 36878 550752
rect 53650 550740 53656 550752
rect 53708 550740 53714 550792
rect 64322 550740 64328 550792
rect 64380 550780 64386 550792
rect 81434 550780 81440 550792
rect 64380 550752 81440 550780
rect 64380 550740 64386 550752
rect 81434 550740 81440 550752
rect 81492 550740 81498 550792
rect 91462 550740 91468 550792
rect 91520 550780 91526 550792
rect 109678 550780 109684 550792
rect 91520 550752 109684 550780
rect 91520 550740 91526 550752
rect 109678 550740 109684 550752
rect 109736 550740 109742 550792
rect 119430 550740 119436 550792
rect 119488 550780 119494 550792
rect 137646 550780 137652 550792
rect 119488 550752 137652 550780
rect 119488 550740 119494 550752
rect 137646 550740 137652 550752
rect 137704 550740 137710 550792
rect 156322 550740 156328 550792
rect 156380 550780 156386 550792
rect 178678 550780 178684 550792
rect 156380 550752 178684 550780
rect 156380 550740 156386 550752
rect 178678 550740 178684 550752
rect 178736 550740 178742 550792
rect 232498 550740 232504 550792
rect 232556 550780 232562 550792
rect 249702 550780 249708 550792
rect 232556 550752 249708 550780
rect 232556 550740 232562 550752
rect 249702 550740 249708 550752
rect 249760 550740 249766 550792
rect 260098 550740 260104 550792
rect 260156 550780 260162 550792
rect 277670 550780 277676 550792
rect 260156 550752 277676 550780
rect 260156 550740 260162 550752
rect 277670 550740 277676 550752
rect 277728 550740 277734 550792
rect 287514 550740 287520 550792
rect 287572 550780 287578 550792
rect 305362 550780 305368 550792
rect 287572 550752 305368 550780
rect 287572 550740 287578 550752
rect 305362 550740 305368 550752
rect 305420 550740 305426 550792
rect 345658 550740 345664 550792
rect 345716 550780 345722 550792
rect 361666 550780 361672 550792
rect 345716 550752 361672 550780
rect 345716 550740 345722 550752
rect 361666 550740 361672 550752
rect 361724 550740 361730 550792
rect 371510 550740 371516 550792
rect 371568 550780 371574 550792
rect 389358 550780 389364 550792
rect 371568 550752 389364 550780
rect 371568 550740 371574 550752
rect 389358 550740 389364 550752
rect 389416 550740 389422 550792
rect 399478 550740 399484 550792
rect 399536 550780 399542 550792
rect 417694 550780 417700 550792
rect 399536 550752 417700 550780
rect 399536 550740 399542 550752
rect 417694 550740 417700 550752
rect 417752 550740 417758 550792
rect 456150 550740 456156 550792
rect 456208 550780 456214 550792
rect 473354 550780 473360 550792
rect 456208 550752 473360 550780
rect 456208 550740 456214 550752
rect 473354 550740 473360 550752
rect 473412 550740 473418 550792
rect 483474 550740 483480 550792
rect 483532 550780 483538 550792
rect 501690 550780 501696 550792
rect 483532 550752 501696 550780
rect 483532 550740 483538 550752
rect 501690 550740 501696 550752
rect 501748 550740 501754 550792
rect 36998 550672 37004 550724
rect 37056 550712 37062 550724
rect 63310 550712 63316 550724
rect 37056 550684 63316 550712
rect 37056 550672 37062 550684
rect 63310 550672 63316 550684
rect 63368 550672 63374 550724
rect 66898 550672 66904 550724
rect 66956 550712 66962 550724
rect 91094 550712 91100 550724
rect 66956 550684 91100 550712
rect 66956 550672 66962 550684
rect 91094 550672 91100 550684
rect 91152 550672 91158 550724
rect 94498 550672 94504 550724
rect 94556 550712 94562 550724
rect 119338 550712 119344 550724
rect 94556 550684 119344 550712
rect 94556 550672 94562 550684
rect 119338 550672 119344 550684
rect 119396 550672 119402 550724
rect 120718 550672 120724 550724
rect 120776 550712 120782 550724
rect 147306 550712 147312 550724
rect 120776 550684 147312 550712
rect 120776 550672 120782 550684
rect 147306 550672 147312 550684
rect 147364 550672 147370 550724
rect 148410 550672 148416 550724
rect 148468 550712 148474 550724
rect 175366 550712 175372 550724
rect 148468 550684 175372 550712
rect 148468 550672 148474 550684
rect 175366 550672 175372 550684
rect 175424 550672 175430 550724
rect 177298 550672 177304 550724
rect 177356 550712 177362 550724
rect 203334 550712 203340 550724
rect 177356 550684 203340 550712
rect 177356 550672 177362 550684
rect 203334 550672 203340 550684
rect 203392 550672 203398 550724
rect 204898 550672 204904 550724
rect 204956 550712 204962 550724
rect 231026 550712 231032 550724
rect 204956 550684 231032 550712
rect 204956 550672 204962 550684
rect 231026 550672 231032 550684
rect 231084 550672 231090 550724
rect 232590 550672 232596 550724
rect 232648 550712 232654 550724
rect 259362 550712 259368 550724
rect 232648 550684 259368 550712
rect 232648 550672 232654 550684
rect 259362 550672 259368 550684
rect 259420 550672 259426 550724
rect 268010 550672 268016 550724
rect 268068 550712 268074 550724
rect 287698 550712 287704 550724
rect 268068 550684 287704 550712
rect 268068 550672 268074 550684
rect 287698 550672 287704 550684
rect 287756 550672 287762 550724
rect 315482 550672 315488 550724
rect 315540 550712 315546 550724
rect 333698 550712 333704 550724
rect 315540 550684 333704 550712
rect 315540 550672 315546 550684
rect 333698 550672 333704 550684
rect 333756 550672 333762 550724
rect 352006 550672 352012 550724
rect 352064 550712 352070 550724
rect 374638 550712 374644 550724
rect 352064 550684 374644 550712
rect 352064 550672 352070 550684
rect 374638 550672 374644 550684
rect 374696 550672 374702 550724
rect 428458 550672 428464 550724
rect 428516 550712 428522 550724
rect 445662 550712 445668 550724
rect 428516 550684 445668 550712
rect 428516 550672 428522 550684
rect 445662 550672 445668 550684
rect 445720 550672 445726 550724
rect 464338 550672 464344 550724
rect 464396 550712 464402 550724
rect 483658 550712 483664 550724
rect 464396 550684 483664 550712
rect 464396 550672 464402 550684
rect 483658 550672 483664 550684
rect 483716 550672 483722 550724
rect 511442 550672 511448 550724
rect 511500 550712 511506 550724
rect 529658 550712 529664 550724
rect 511500 550684 529664 550712
rect 511500 550672 511506 550684
rect 529658 550672 529664 550684
rect 529716 550672 529722 550724
rect 542998 550672 543004 550724
rect 543056 550712 543062 550724
rect 557534 550712 557540 550724
rect 543056 550684 557540 550712
rect 543056 550672 543062 550684
rect 557534 550672 557540 550684
rect 557592 550672 557598 550724
rect 212350 550604 212356 550656
rect 212408 550644 212414 550656
rect 232682 550644 232688 550656
rect 212408 550616 232688 550644
rect 212408 550604 212414 550616
rect 232682 550604 232688 550616
rect 232740 550604 232746 550656
rect 260190 550604 260196 550656
rect 260248 550644 260254 550656
rect 287330 550644 287336 550656
rect 260248 550616 287336 550644
rect 260248 550604 260254 550616
rect 287330 550604 287336 550616
rect 287388 550604 287394 550656
rect 289078 550604 289084 550656
rect 289136 550644 289142 550656
rect 315022 550644 315028 550656
rect 289136 550616 315028 550644
rect 289136 550604 289142 550616
rect 315022 550604 315028 550616
rect 315080 550604 315086 550656
rect 316678 550604 316684 550656
rect 316736 550644 316742 550656
rect 343358 550644 343364 550656
rect 316736 550616 343364 550644
rect 316736 550604 316742 550616
rect 343358 550604 343364 550616
rect 343416 550604 343422 550656
rect 344278 550604 344284 550656
rect 344336 550644 344342 550656
rect 371326 550644 371332 550656
rect 344336 550616 371332 550644
rect 344336 550604 344342 550616
rect 371326 550604 371332 550616
rect 371384 550604 371390 550656
rect 373258 550604 373264 550656
rect 373316 550644 373322 550656
rect 399018 550644 399024 550656
rect 373316 550616 399024 550644
rect 373316 550604 373322 550616
rect 399018 550604 399024 550616
rect 399076 550604 399082 550656
rect 400858 550604 400864 550656
rect 400916 550644 400922 550656
rect 427354 550644 427360 550656
rect 400916 550616 427360 550644
rect 400916 550604 400922 550616
rect 427354 550604 427360 550616
rect 427412 550604 427418 550656
rect 428550 550604 428556 550656
rect 428608 550644 428614 550656
rect 455322 550644 455328 550656
rect 428608 550616 455328 550644
rect 428608 550604 428614 550616
rect 455322 550604 455328 550616
rect 455380 550604 455386 550656
rect 456058 550604 456064 550656
rect 456116 550644 456122 550656
rect 483014 550644 483020 550656
rect 456116 550616 483020 550644
rect 456116 550604 456122 550616
rect 483014 550604 483020 550616
rect 483072 550604 483078 550656
rect 485038 550604 485044 550656
rect 485096 550644 485102 550656
rect 511350 550644 511356 550656
rect 485096 550616 511356 550644
rect 485096 550604 485102 550616
rect 511350 550604 511356 550616
rect 511408 550604 511414 550656
rect 512638 550604 512644 550656
rect 512696 550644 512702 550656
rect 539318 550644 539324 550656
rect 512696 550616 539324 550644
rect 512696 550604 512702 550616
rect 539318 550604 539324 550616
rect 539376 550604 539382 550656
rect 540238 550604 540244 550656
rect 540296 550644 540302 550656
rect 567194 550644 567200 550656
rect 540296 550616 567200 550644
rect 540296 550604 540302 550616
rect 567194 550604 567200 550616
rect 567252 550604 567258 550656
rect 37918 548496 37924 548548
rect 37976 548536 37982 548548
rect 545758 548536 545764 548548
rect 37976 548508 545764 548536
rect 37976 548496 37982 548508
rect 545758 548496 545764 548508
rect 545816 548496 545822 548548
rect 35618 547884 35624 547936
rect 35676 547924 35682 547936
rect 36906 547924 36912 547936
rect 35676 547896 36912 547924
rect 35676 547884 35682 547896
rect 36906 547884 36912 547896
rect 36964 547884 36970 547936
rect 63586 533604 63592 533656
rect 63644 533644 63650 533656
rect 64322 533644 64328 533656
rect 63644 533616 64328 533644
rect 63644 533604 63650 533616
rect 64322 533604 64328 533616
rect 64380 533604 64386 533656
rect 455690 533604 455696 533656
rect 455748 533644 455754 533656
rect 456150 533644 456156 533656
rect 455748 533616 456156 533644
rect 455748 533604 455754 533616
rect 456150 533604 456156 533616
rect 456208 533604 456214 533656
rect 316770 530680 316776 530732
rect 316828 530720 316834 530732
rect 323670 530720 323676 530732
rect 316828 530692 323676 530720
rect 316828 530680 316834 530692
rect 323670 530680 323676 530692
rect 323728 530680 323734 530732
rect 428642 530544 428648 530596
rect 428700 530584 428706 530596
rect 435726 530584 435732 530596
rect 428700 530556 435732 530584
rect 428700 530544 428706 530556
rect 435726 530544 435732 530556
rect 435784 530544 435790 530596
rect 287698 530272 287704 530324
rect 287756 530312 287762 530324
rect 295702 530312 295708 530324
rect 287756 530284 295708 530312
rect 287756 530272 287762 530284
rect 295702 530272 295708 530284
rect 295760 530272 295766 530324
rect 232682 530204 232688 530256
rect 232740 530244 232746 530256
rect 239766 530244 239772 530256
rect 232740 530216 239772 530244
rect 232740 530204 232746 530216
rect 239766 530204 239772 530216
rect 239824 530204 239830 530256
rect 512730 530204 512736 530256
rect 512788 530244 512794 530256
rect 519630 530244 519636 530256
rect 512788 530216 519636 530244
rect 512788 530204 512794 530216
rect 519630 530204 519636 530216
rect 519688 530204 519694 530256
rect 483658 530136 483664 530188
rect 483716 530176 483722 530188
rect 491662 530176 491668 530188
rect 483716 530148 491668 530176
rect 483716 530136 483722 530148
rect 491662 530136 491668 530148
rect 491720 530136 491726 530188
rect 13722 529864 13728 529916
rect 13780 529904 13786 529916
rect 66254 529904 66260 529916
rect 13780 529876 66260 529904
rect 13780 529864 13786 529876
rect 66254 529864 66260 529876
rect 66312 529864 66318 529916
rect 97902 529864 97908 529916
rect 97960 529904 97966 529916
rect 149054 529904 149060 529916
rect 97960 529876 149060 529904
rect 97960 529864 97966 529876
rect 149054 529864 149060 529876
rect 149112 529864 149118 529916
rect 154482 529864 154488 529916
rect 154540 529904 154546 529916
rect 205634 529904 205640 529916
rect 154540 529876 205640 529904
rect 154540 529864 154546 529876
rect 205634 529864 205640 529876
rect 205692 529864 205698 529916
rect 209682 529864 209688 529916
rect 209740 529904 209746 529916
rect 262214 529904 262220 529916
rect 209740 529876 262220 529904
rect 209740 529864 209746 529876
rect 262214 529864 262220 529876
rect 262272 529864 262278 529916
rect 266262 529864 266268 529916
rect 266320 529904 266326 529916
rect 317414 529904 317420 529916
rect 266320 529876 317420 529904
rect 266320 529864 266326 529876
rect 317414 529864 317420 529876
rect 317472 529864 317478 529916
rect 322842 529864 322848 529916
rect 322900 529904 322906 529916
rect 373994 529904 374000 529916
rect 322900 529876 374000 529904
rect 322900 529864 322906 529876
rect 373994 529864 374000 529876
rect 374052 529864 374058 529916
rect 405642 529864 405648 529916
rect 405700 529904 405706 529916
rect 458174 529904 458180 529916
rect 405700 529876 458180 529904
rect 405700 529864 405706 529876
rect 458174 529864 458180 529876
rect 458232 529864 458238 529916
rect 489822 529864 489828 529916
rect 489880 529904 489886 529916
rect 542354 529904 542360 529916
rect 489880 529876 542360 529904
rect 489880 529864 489886 529876
rect 542354 529864 542360 529876
rect 542412 529864 542418 529916
rect 35618 529796 35624 529848
rect 35676 529836 35682 529848
rect 36814 529836 36820 529848
rect 35676 529808 36820 529836
rect 35676 529796 35682 529808
rect 36814 529796 36820 529808
rect 36872 529796 36878 529848
rect 42702 529796 42708 529848
rect 42760 529836 42766 529848
rect 93854 529836 93860 529848
rect 42760 529808 93860 529836
rect 42760 529796 42766 529808
rect 93854 529796 93860 529808
rect 93912 529796 93918 529848
rect 126882 529796 126888 529848
rect 126940 529836 126946 529848
rect 178034 529836 178040 529848
rect 126940 529808 178040 529836
rect 126940 529796 126946 529808
rect 178034 529796 178040 529808
rect 178092 529796 178098 529848
rect 182082 529796 182088 529848
rect 182140 529836 182146 529848
rect 233234 529836 233240 529848
rect 182140 529808 233240 529836
rect 182140 529796 182146 529808
rect 233234 529796 233240 529808
rect 233292 529796 233298 529848
rect 238662 529796 238668 529848
rect 238720 529836 238726 529848
rect 289814 529836 289820 529848
rect 238720 529808 289820 529836
rect 238720 529796 238726 529808
rect 289814 529796 289820 529808
rect 289872 529796 289878 529848
rect 293862 529796 293868 529848
rect 293920 529836 293926 529848
rect 293920 529808 335354 529836
rect 293920 529796 293926 529808
rect 70302 529728 70308 529780
rect 70360 529768 70366 529780
rect 121454 529768 121460 529780
rect 70360 529740 121460 529768
rect 70360 529728 70366 529740
rect 121454 529728 121460 529740
rect 121512 529728 121518 529780
rect 335326 529768 335354 529808
rect 343542 529796 343548 529848
rect 343600 529836 343606 529848
rect 345658 529836 345664 529848
rect 343600 529808 345664 529836
rect 343600 529796 343606 529808
rect 345658 529796 345664 529808
rect 345716 529796 345722 529848
rect 350442 529796 350448 529848
rect 350500 529836 350506 529848
rect 401594 529836 401600 529848
rect 350500 529808 401600 529836
rect 350500 529796 350506 529808
rect 401594 529796 401600 529808
rect 401652 529796 401658 529848
rect 434622 529796 434628 529848
rect 434680 529836 434686 529848
rect 485774 529836 485780 529848
rect 434680 529808 485780 529836
rect 434680 529796 434686 529808
rect 485774 529796 485780 529808
rect 485832 529796 485838 529848
rect 518802 529796 518808 529848
rect 518860 529836 518866 529848
rect 569954 529836 569960 529848
rect 518860 529808 569960 529836
rect 518860 529796 518866 529808
rect 569954 529796 569960 529808
rect 570012 529796 570018 529848
rect 345014 529768 345020 529780
rect 335326 529740 345020 529768
rect 345014 529728 345020 529740
rect 345072 529728 345078 529780
rect 378042 529728 378048 529780
rect 378100 529768 378106 529780
rect 429194 529768 429200 529780
rect 378100 529740 429200 529768
rect 378100 529728 378106 529740
rect 429194 529728 429200 529740
rect 429252 529728 429258 529780
rect 462222 529728 462228 529780
rect 462280 529768 462286 529780
rect 513374 529768 513380 529780
rect 462280 529740 513380 529768
rect 462280 529728 462286 529740
rect 513374 529728 513380 529740
rect 513432 529728 513438 529780
rect 178678 527076 178684 527128
rect 178736 527116 178742 527128
rect 184014 527116 184020 527128
rect 178736 527088 184020 527116
rect 178736 527076 178742 527088
rect 184014 527076 184020 527088
rect 184072 527076 184078 527128
rect 374638 527076 374644 527128
rect 374696 527116 374702 527128
rect 379698 527116 379704 527128
rect 374696 527088 379704 527116
rect 374696 527076 374702 527088
rect 379698 527076 379704 527088
rect 379756 527076 379762 527128
rect 539318 527076 539324 527128
rect 539376 527116 539382 527128
rect 542998 527116 543004 527128
rect 539376 527088 543004 527116
rect 539376 527076 539382 527088
rect 542998 527076 543004 527088
rect 543056 527076 543062 527128
rect 15194 527008 15200 527060
rect 15252 527048 15258 527060
rect 43990 527048 43996 527060
rect 15252 527020 43996 527048
rect 15252 527008 15258 527020
rect 43990 527008 43996 527020
rect 44048 527008 44054 527060
rect 71038 527008 71044 527060
rect 71096 527048 71102 527060
rect 567194 527048 567200 527060
rect 71096 527020 567200 527048
rect 71096 527008 71102 527020
rect 567194 527008 567200 527020
rect 567252 527008 567258 527060
rect 25682 526940 25688 526992
rect 25740 526980 25746 526992
rect 36998 526980 37004 526992
rect 25740 526952 37004 526980
rect 25740 526940 25746 526952
rect 36998 526940 37004 526952
rect 37056 526940 37062 526992
rect 53650 526940 53656 526992
rect 53708 526980 53714 526992
rect 66898 526980 66904 526992
rect 53708 526952 66904 526980
rect 53708 526940 53714 526952
rect 66898 526940 66904 526952
rect 66956 526940 66962 526992
rect 71866 526940 71872 526992
rect 71924 526980 71930 526992
rect 100018 526980 100024 526992
rect 71924 526952 100024 526980
rect 71924 526940 71930 526952
rect 100018 526940 100024 526952
rect 100076 526940 100082 526992
rect 127986 526980 127992 526992
rect 103486 526952 127992 526980
rect 42886 526872 42892 526924
rect 42944 526912 42950 526924
rect 71958 526912 71964 526924
rect 42944 526884 71964 526912
rect 42944 526872 42950 526884
rect 71958 526872 71964 526884
rect 72016 526872 72022 526924
rect 81986 526872 81992 526924
rect 82044 526912 82050 526924
rect 94498 526912 94504 526924
rect 82044 526884 94504 526912
rect 82044 526872 82050 526884
rect 94498 526872 94504 526884
rect 94556 526872 94562 526924
rect 99466 526872 99472 526924
rect 99524 526912 99530 526924
rect 103486 526912 103514 526952
rect 127986 526940 127992 526952
rect 128044 526940 128050 526992
rect 155954 526980 155960 526992
rect 132466 526952 155960 526980
rect 99524 526884 103514 526912
rect 99524 526872 99530 526884
rect 109678 526872 109684 526924
rect 109736 526912 109742 526924
rect 120718 526912 120724 526924
rect 109736 526884 120724 526912
rect 109736 526872 109742 526884
rect 120718 526872 120724 526884
rect 120776 526872 120782 526924
rect 127066 526872 127072 526924
rect 127124 526912 127130 526924
rect 132466 526912 132494 526952
rect 155954 526940 155960 526952
rect 156012 526940 156018 526992
rect 165982 526940 165988 526992
rect 166040 526980 166046 526992
rect 177298 526980 177304 526992
rect 166040 526952 177304 526980
rect 166040 526940 166046 526952
rect 177298 526940 177304 526952
rect 177356 526940 177362 526992
rect 183646 526940 183652 526992
rect 183704 526980 183710 526992
rect 211706 526980 211712 526992
rect 183704 526952 211712 526980
rect 183704 526940 183710 526952
rect 211706 526940 211712 526952
rect 211764 526940 211770 526992
rect 221918 526940 221924 526992
rect 221976 526980 221982 526992
rect 232590 526980 232596 526992
rect 221976 526952 232596 526980
rect 221976 526940 221982 526952
rect 232590 526940 232596 526952
rect 232648 526940 232654 526992
rect 238846 526940 238852 526992
rect 238904 526980 238910 526992
rect 268010 526980 268016 526992
rect 238904 526952 268016 526980
rect 238904 526940 238910 526952
rect 268010 526940 268016 526952
rect 268068 526940 268074 526992
rect 277670 526940 277676 526992
rect 277728 526980 277734 526992
rect 289078 526980 289084 526992
rect 277728 526952 289084 526980
rect 277728 526940 277734 526952
rect 289078 526940 289084 526952
rect 289136 526940 289142 526992
rect 306006 526940 306012 526992
rect 306064 526980 306070 526992
rect 316678 526980 316684 526992
rect 306064 526952 316684 526980
rect 306064 526940 306070 526952
rect 316678 526940 316684 526952
rect 316736 526940 316742 526992
rect 323026 526940 323032 526992
rect 323084 526980 323090 526992
rect 352006 526980 352012 526992
rect 323084 526952 352012 526980
rect 323084 526940 323090 526952
rect 352006 526940 352012 526952
rect 352064 526940 352070 526992
rect 361666 526940 361672 526992
rect 361724 526980 361730 526992
rect 373258 526980 373264 526992
rect 361724 526952 373264 526980
rect 361724 526940 361730 526952
rect 373258 526940 373264 526952
rect 373316 526940 373322 526992
rect 379606 526940 379612 526992
rect 379664 526980 379670 526992
rect 408034 526980 408040 526992
rect 379664 526952 408040 526980
rect 379664 526940 379670 526952
rect 408034 526940 408040 526952
rect 408092 526940 408098 526992
rect 417694 526940 417700 526992
rect 417752 526980 417758 526992
rect 428550 526980 428556 526992
rect 417752 526952 428556 526980
rect 417752 526940 417758 526952
rect 428550 526940 428556 526952
rect 428608 526940 428614 526992
rect 434806 526940 434812 526992
rect 434864 526980 434870 526992
rect 463786 526980 463792 526992
rect 434864 526952 463792 526980
rect 434864 526940 434870 526952
rect 463786 526940 463792 526952
rect 463844 526940 463850 526992
rect 473998 526940 474004 526992
rect 474056 526980 474062 526992
rect 485038 526980 485044 526992
rect 474056 526952 485044 526980
rect 474056 526940 474062 526952
rect 485038 526940 485044 526952
rect 485096 526940 485102 526992
rect 501690 526940 501696 526992
rect 501748 526980 501754 526992
rect 512638 526980 512644 526992
rect 501748 526952 512644 526980
rect 501748 526940 501754 526952
rect 512638 526940 512644 526952
rect 512696 526940 512702 526992
rect 518986 526940 518992 526992
rect 519044 526980 519050 526992
rect 547874 526980 547880 526992
rect 519044 526952 547880 526980
rect 519044 526940 519050 526952
rect 547874 526940 547880 526952
rect 547932 526940 547938 526992
rect 127124 526884 132494 526912
rect 127124 526872 127130 526884
rect 137646 526872 137652 526924
rect 137704 526912 137710 526924
rect 148410 526912 148416 526924
rect 137704 526884 148416 526912
rect 137704 526872 137710 526884
rect 148410 526872 148416 526884
rect 148468 526872 148474 526924
rect 193674 526872 193680 526924
rect 193732 526912 193738 526924
rect 204898 526912 204904 526924
rect 193732 526884 204904 526912
rect 193732 526872 193738 526884
rect 204898 526872 204904 526884
rect 204956 526872 204962 526924
rect 249702 526872 249708 526924
rect 249760 526912 249766 526924
rect 260190 526912 260196 526924
rect 249760 526884 260196 526912
rect 249760 526872 249766 526884
rect 260190 526872 260196 526884
rect 260248 526872 260254 526924
rect 333698 526872 333704 526924
rect 333756 526912 333762 526924
rect 344278 526912 344284 526924
rect 333756 526884 344284 526912
rect 333756 526872 333762 526884
rect 344278 526872 344284 526884
rect 344336 526872 344342 526924
rect 390002 526872 390008 526924
rect 390060 526912 390066 526924
rect 400858 526912 400864 526924
rect 390060 526884 400864 526912
rect 390060 526872 390066 526884
rect 400858 526872 400864 526884
rect 400916 526872 400922 526924
rect 445662 526872 445668 526924
rect 445720 526912 445726 526924
rect 456058 526912 456064 526924
rect 445720 526884 456064 526912
rect 445720 526872 445726 526884
rect 456058 526872 456064 526884
rect 456116 526872 456122 526924
rect 529658 526872 529664 526924
rect 529716 526912 529722 526924
rect 540238 526912 540244 526924
rect 529716 526884 540244 526912
rect 529716 526872 529722 526884
rect 540238 526872 540244 526884
rect 540296 526872 540302 526924
rect 36722 526804 36728 526856
rect 36780 526844 36786 526856
rect 557534 526844 557540 526856
rect 36780 526816 557540 526844
rect 36780 526804 36786 526816
rect 557534 526804 557540 526816
rect 557592 526804 557598 526856
rect 16022 523676 16028 523728
rect 16080 523716 16086 523728
rect 547874 523716 547880 523728
rect 16080 523688 547880 523716
rect 16080 523676 16086 523688
rect 547874 523676 547880 523688
rect 547932 523676 547938 523728
rect 25682 523200 25688 523252
rect 25740 523240 25746 523252
rect 71038 523240 71044 523252
rect 25740 523212 71044 523240
rect 25740 523200 25746 523212
rect 71038 523200 71044 523212
rect 71096 523200 71102 523252
rect 212350 523200 212356 523252
rect 212408 523240 212414 523252
rect 232682 523240 232688 523252
rect 212408 523212 232688 523240
rect 212408 523200 212414 523212
rect 232682 523200 232688 523212
rect 232740 523200 232746 523252
rect 296346 523200 296352 523252
rect 296404 523240 296410 523252
rect 316770 523240 316776 523252
rect 296404 523212 316776 523240
rect 296404 523200 296410 523212
rect 316770 523200 316776 523212
rect 316828 523200 316834 523252
rect 408034 523200 408040 523252
rect 408092 523240 408098 523252
rect 428642 523240 428648 523252
rect 408092 523212 428648 523240
rect 408092 523200 408098 523212
rect 428642 523200 428648 523212
rect 428700 523200 428706 523252
rect 492030 523200 492036 523252
rect 492088 523240 492094 523252
rect 512730 523240 512736 523252
rect 492088 523212 512736 523240
rect 492088 523200 492094 523212
rect 512730 523200 512736 523212
rect 512788 523200 512794 523252
rect 36722 523132 36728 523184
rect 36780 523172 36786 523184
rect 53650 523172 53656 523184
rect 36780 523144 53656 523172
rect 36780 523132 36786 523144
rect 53650 523132 53656 523144
rect 53708 523132 53714 523184
rect 148410 523132 148416 523184
rect 148468 523172 148474 523184
rect 165706 523172 165712 523184
rect 148468 523144 165712 523172
rect 148468 523132 148474 523144
rect 165706 523132 165712 523144
rect 165764 523132 165770 523184
rect 175458 523132 175464 523184
rect 175516 523172 175522 523184
rect 193674 523172 193680 523184
rect 175516 523144 193680 523172
rect 175516 523132 175522 523144
rect 193674 523132 193680 523144
rect 193732 523132 193738 523184
rect 203518 523132 203524 523184
rect 203576 523172 203582 523184
rect 221366 523172 221372 523184
rect 203576 523144 221372 523172
rect 203576 523132 203582 523144
rect 221366 523132 221372 523144
rect 221424 523132 221430 523184
rect 260190 523132 260196 523184
rect 260248 523172 260254 523184
rect 277670 523172 277676 523184
rect 260248 523144 277676 523172
rect 260248 523132 260254 523144
rect 277670 523132 277676 523144
rect 277728 523132 277734 523184
rect 287514 523132 287520 523184
rect 287572 523172 287578 523184
rect 305362 523172 305368 523184
rect 287572 523144 305368 523172
rect 287572 523132 287578 523144
rect 305362 523132 305368 523144
rect 305420 523132 305426 523184
rect 345658 523132 345664 523184
rect 345716 523172 345722 523184
rect 361666 523172 361672 523184
rect 345716 523144 361672 523172
rect 345716 523132 345722 523144
rect 361666 523132 361672 523144
rect 361724 523132 361730 523184
rect 371510 523132 371516 523184
rect 371568 523172 371574 523184
rect 389358 523172 389364 523184
rect 371568 523144 389364 523172
rect 371568 523132 371574 523144
rect 389358 523132 389364 523144
rect 389416 523132 389422 523184
rect 399478 523132 399484 523184
rect 399536 523172 399542 523184
rect 417694 523172 417700 523184
rect 399536 523144 417700 523172
rect 399536 523132 399542 523144
rect 417694 523132 417700 523144
rect 417752 523132 417758 523184
rect 456150 523132 456156 523184
rect 456208 523172 456214 523184
rect 473354 523172 473360 523184
rect 456208 523144 473360 523172
rect 456208 523132 456214 523144
rect 473354 523132 473360 523144
rect 473412 523132 473418 523184
rect 483474 523132 483480 523184
rect 483532 523172 483538 523184
rect 501690 523172 501696 523184
rect 483532 523144 501696 523172
rect 483532 523132 483538 523144
rect 501690 523132 501696 523144
rect 501748 523132 501754 523184
rect 36998 523064 37004 523116
rect 37056 523104 37062 523116
rect 63310 523104 63316 523116
rect 37056 523076 63316 523104
rect 37056 523064 37062 523076
rect 63310 523064 63316 523076
rect 63368 523064 63374 523116
rect 64322 523064 64328 523116
rect 64380 523104 64386 523116
rect 81434 523104 81440 523116
rect 64380 523076 81440 523104
rect 64380 523064 64386 523076
rect 81434 523064 81440 523076
rect 81492 523064 81498 523116
rect 91462 523064 91468 523116
rect 91520 523104 91526 523116
rect 109678 523104 109684 523116
rect 91520 523076 109684 523104
rect 91520 523064 91526 523076
rect 109678 523064 109684 523076
rect 109736 523064 109742 523116
rect 119430 523064 119436 523116
rect 119488 523104 119494 523116
rect 137646 523104 137652 523116
rect 119488 523076 137652 523104
rect 119488 523064 119494 523076
rect 137646 523064 137652 523076
rect 137704 523064 137710 523116
rect 156322 523064 156328 523116
rect 156380 523104 156386 523116
rect 178678 523104 178684 523116
rect 156380 523076 178684 523104
rect 156380 523064 156386 523076
rect 178678 523064 178684 523076
rect 178736 523064 178742 523116
rect 232498 523064 232504 523116
rect 232556 523104 232562 523116
rect 249702 523104 249708 523116
rect 232556 523076 249708 523104
rect 232556 523064 232562 523076
rect 249702 523064 249708 523076
rect 249760 523064 249766 523116
rect 268010 523064 268016 523116
rect 268068 523104 268074 523116
rect 287698 523104 287704 523116
rect 268068 523076 287704 523104
rect 268068 523064 268074 523076
rect 287698 523064 287704 523076
rect 287756 523064 287762 523116
rect 315482 523064 315488 523116
rect 315540 523104 315546 523116
rect 333698 523104 333704 523116
rect 315540 523076 333704 523104
rect 315540 523064 315546 523076
rect 333698 523064 333704 523076
rect 333756 523064 333762 523116
rect 352006 523064 352012 523116
rect 352064 523104 352070 523116
rect 374638 523104 374644 523116
rect 352064 523076 374644 523104
rect 352064 523064 352070 523076
rect 374638 523064 374644 523076
rect 374696 523064 374702 523116
rect 428550 523064 428556 523116
rect 428608 523104 428614 523116
rect 445662 523104 445668 523116
rect 428608 523076 445668 523104
rect 428608 523064 428614 523076
rect 445662 523064 445668 523076
rect 445720 523064 445726 523116
rect 464338 523064 464344 523116
rect 464396 523104 464402 523116
rect 483658 523104 483664 523116
rect 464396 523076 483664 523104
rect 464396 523064 464402 523076
rect 483658 523064 483664 523076
rect 483716 523064 483722 523116
rect 511442 523064 511448 523116
rect 511500 523104 511506 523116
rect 529658 523104 529664 523116
rect 511500 523076 529664 523104
rect 511500 523064 511506 523076
rect 529658 523064 529664 523076
rect 529716 523064 529722 523116
rect 542998 523064 543004 523116
rect 543056 523104 543062 523116
rect 557534 523104 557540 523116
rect 543056 523076 557540 523104
rect 543056 523064 543062 523076
rect 557534 523064 557540 523076
rect 557592 523064 557598 523116
rect 69658 522996 69664 523048
rect 69716 523036 69722 523048
rect 91094 523036 91100 523048
rect 69716 523008 91100 523036
rect 69716 522996 69722 523008
rect 91094 522996 91100 523008
rect 91152 522996 91158 523048
rect 94498 522996 94504 523048
rect 94556 523036 94562 523048
rect 119338 523036 119344 523048
rect 94556 523008 119344 523036
rect 94556 522996 94562 523008
rect 119338 522996 119344 523008
rect 119396 522996 119402 523048
rect 120718 522996 120724 523048
rect 120776 523036 120782 523048
rect 147306 523036 147312 523048
rect 120776 523008 147312 523036
rect 120776 522996 120782 523008
rect 147306 522996 147312 523008
rect 147364 522996 147370 523048
rect 148318 522996 148324 523048
rect 148376 523036 148382 523048
rect 175366 523036 175372 523048
rect 148376 523008 175372 523036
rect 148376 522996 148382 523008
rect 175366 522996 175372 523008
rect 175424 522996 175430 523048
rect 177298 522996 177304 523048
rect 177356 523036 177362 523048
rect 203334 523036 203340 523048
rect 177356 523008 203340 523036
rect 177356 522996 177362 523008
rect 203334 522996 203340 523008
rect 203392 522996 203398 523048
rect 204898 522996 204904 523048
rect 204956 523036 204962 523048
rect 231026 523036 231032 523048
rect 204956 523008 231032 523036
rect 204956 522996 204962 523008
rect 231026 522996 231032 523008
rect 231084 522996 231090 523048
rect 232590 522996 232596 523048
rect 232648 523036 232654 523048
rect 259362 523036 259368 523048
rect 232648 523008 259368 523036
rect 232648 522996 232654 523008
rect 259362 522996 259368 523008
rect 259420 522996 259426 523048
rect 260098 522996 260104 523048
rect 260156 523036 260162 523048
rect 287330 523036 287336 523048
rect 260156 523008 287336 523036
rect 260156 522996 260162 523008
rect 287330 522996 287336 523008
rect 287388 522996 287394 523048
rect 289078 522996 289084 523048
rect 289136 523036 289142 523048
rect 315022 523036 315028 523048
rect 289136 523008 315028 523036
rect 289136 522996 289142 523008
rect 315022 522996 315028 523008
rect 315080 522996 315086 523048
rect 316678 522996 316684 523048
rect 316736 523036 316742 523048
rect 343358 523036 343364 523048
rect 316736 523008 343364 523036
rect 316736 522996 316742 523008
rect 343358 522996 343364 523008
rect 343416 522996 343422 523048
rect 344278 522996 344284 523048
rect 344336 523036 344342 523048
rect 371326 523036 371332 523048
rect 344336 523008 371332 523036
rect 344336 522996 344342 523008
rect 371326 522996 371332 523008
rect 371384 522996 371390 523048
rect 373258 522996 373264 523048
rect 373316 523036 373322 523048
rect 399018 523036 399024 523048
rect 373316 523008 399024 523036
rect 373316 522996 373322 523008
rect 399018 522996 399024 523008
rect 399076 522996 399082 523048
rect 400858 522996 400864 523048
rect 400916 523036 400922 523048
rect 427354 523036 427360 523048
rect 400916 523008 427360 523036
rect 400916 522996 400922 523008
rect 427354 522996 427360 523008
rect 427412 522996 427418 523048
rect 428458 522996 428464 523048
rect 428516 523036 428522 523048
rect 455322 523036 455328 523048
rect 428516 523008 455328 523036
rect 428516 522996 428522 523008
rect 455322 522996 455328 523008
rect 455380 522996 455386 523048
rect 456058 522996 456064 523048
rect 456116 523036 456122 523048
rect 483014 523036 483020 523048
rect 456116 523008 483020 523036
rect 456116 522996 456122 523008
rect 483014 522996 483020 523008
rect 483072 522996 483078 523048
rect 485038 522996 485044 523048
rect 485096 523036 485102 523048
rect 511350 523036 511356 523048
rect 485096 523008 511356 523036
rect 485096 522996 485102 523008
rect 511350 522996 511356 523008
rect 511408 522996 511414 523048
rect 512638 522996 512644 523048
rect 512696 523036 512702 523048
rect 539318 523036 539324 523048
rect 512696 523008 539324 523036
rect 512696 522996 512702 523008
rect 539318 522996 539324 523008
rect 539376 522996 539382 523048
rect 540238 522996 540244 523048
rect 540296 523036 540302 523048
rect 567194 523036 567200 523048
rect 540296 523008 567200 523036
rect 540296 522996 540302 523008
rect 567194 522996 567200 523008
rect 567252 522996 567258 523048
rect 37918 522248 37924 522300
rect 37976 522288 37982 522300
rect 545758 522288 545764 522300
rect 37976 522260 545764 522288
rect 37976 522248 37982 522260
rect 545758 522248 545764 522260
rect 545816 522248 545822 522300
rect 35618 521704 35624 521756
rect 35676 521744 35682 521756
rect 36814 521744 36820 521756
rect 35676 521716 36820 521744
rect 35676 521704 35682 521716
rect 36814 521704 36820 521716
rect 36872 521704 36878 521756
rect 42702 520344 42708 520396
rect 42760 520384 42766 520396
rect 93854 520384 93860 520396
rect 42760 520356 93860 520384
rect 42760 520344 42766 520356
rect 93854 520344 93860 520356
rect 93912 520344 93918 520396
rect 155862 520344 155868 520396
rect 155920 520384 155926 520396
rect 205634 520384 205640 520396
rect 155920 520356 205640 520384
rect 155920 520344 155926 520356
rect 205634 520344 205640 520356
rect 205692 520344 205698 520396
rect 238662 520344 238668 520396
rect 238720 520384 238726 520396
rect 289814 520384 289820 520396
rect 238720 520356 289820 520384
rect 238720 520344 238726 520356
rect 289814 520344 289820 520356
rect 289872 520344 289878 520396
rect 322842 520344 322848 520396
rect 322900 520384 322906 520396
rect 373994 520384 374000 520396
rect 322900 520356 374000 520384
rect 322900 520344 322906 520356
rect 373994 520344 374000 520356
rect 374052 520344 374058 520396
rect 434622 520344 434628 520396
rect 434680 520384 434686 520396
rect 485774 520384 485780 520396
rect 434680 520356 485780 520384
rect 434680 520344 434686 520356
rect 485774 520344 485780 520356
rect 485832 520344 485838 520396
rect 13722 520276 13728 520328
rect 13780 520316 13786 520328
rect 66254 520316 66260 520328
rect 13780 520288 66260 520316
rect 13780 520276 13786 520288
rect 66254 520276 66260 520288
rect 66312 520276 66318 520328
rect 70302 520276 70308 520328
rect 70360 520316 70366 520328
rect 121454 520316 121460 520328
rect 70360 520288 121460 520316
rect 70360 520276 70366 520288
rect 121454 520276 121460 520288
rect 121512 520276 121518 520328
rect 126882 520276 126888 520328
rect 126940 520316 126946 520328
rect 178034 520316 178040 520328
rect 126940 520288 178040 520316
rect 126940 520276 126946 520288
rect 178034 520276 178040 520288
rect 178092 520276 178098 520328
rect 209682 520276 209688 520328
rect 209740 520316 209746 520328
rect 262214 520316 262220 520328
rect 209740 520288 262220 520316
rect 209740 520276 209746 520288
rect 262214 520276 262220 520288
rect 262272 520276 262278 520328
rect 293862 520276 293868 520328
rect 293920 520316 293926 520328
rect 345014 520316 345020 520328
rect 293920 520288 345020 520316
rect 293920 520276 293926 520288
rect 345014 520276 345020 520288
rect 345072 520276 345078 520328
rect 350442 520276 350448 520328
rect 350500 520316 350506 520328
rect 401594 520316 401600 520328
rect 350500 520288 401600 520316
rect 350500 520276 350506 520288
rect 401594 520276 401600 520288
rect 401652 520276 401658 520328
rect 407850 520276 407856 520328
rect 407908 520316 407914 520328
rect 458174 520316 458180 520328
rect 407908 520288 458180 520316
rect 407908 520276 407914 520288
rect 458174 520276 458180 520288
rect 458232 520276 458238 520328
rect 518802 520276 518808 520328
rect 518860 520316 518866 520328
rect 569954 520316 569960 520328
rect 518860 520288 569960 520316
rect 518860 520276 518866 520288
rect 569954 520276 569960 520288
rect 570012 520276 570018 520328
rect 154482 518848 154488 518900
rect 154540 518888 154546 518900
rect 155862 518888 155868 518900
rect 154540 518860 155868 518888
rect 154540 518848 154546 518860
rect 155862 518848 155868 518860
rect 155920 518848 155926 518900
rect 540882 509192 540888 509244
rect 540940 509232 540946 509244
rect 542354 509232 542360 509244
rect 540940 509204 542360 509232
rect 540940 509192 540946 509204
rect 542354 509192 542360 509204
rect 542412 509192 542418 509244
rect 63586 505588 63592 505640
rect 63644 505628 63650 505640
rect 64322 505628 64328 505640
rect 63644 505600 64328 505628
rect 63644 505588 63650 505600
rect 64322 505588 64328 505600
rect 64380 505588 64386 505640
rect 147674 505588 147680 505640
rect 147732 505628 147738 505640
rect 148410 505628 148416 505640
rect 147732 505600 148416 505628
rect 147732 505588 147738 505600
rect 148410 505588 148416 505600
rect 148468 505588 148474 505640
rect 259730 505588 259736 505640
rect 259788 505628 259794 505640
rect 260190 505628 260196 505640
rect 259788 505600 260196 505628
rect 259788 505588 259794 505600
rect 260190 505588 260196 505600
rect 260248 505588 260254 505640
rect 455690 505588 455696 505640
rect 455748 505628 455754 505640
rect 456150 505628 456156 505640
rect 455748 505600 456156 505628
rect 455748 505588 455754 505600
rect 456150 505588 456156 505600
rect 456208 505588 456214 505640
rect 287698 504568 287704 504620
rect 287756 504608 287762 504620
rect 295702 504608 295708 504620
rect 287756 504580 295708 504608
rect 287756 504568 287762 504580
rect 295702 504568 295708 504580
rect 295760 504568 295766 504620
rect 428642 504364 428648 504416
rect 428700 504404 428706 504416
rect 435726 504404 435732 504416
rect 428700 504376 435732 504404
rect 428700 504364 428706 504376
rect 435726 504364 435732 504376
rect 435784 504364 435790 504416
rect 483658 504296 483664 504348
rect 483716 504336 483722 504348
rect 491662 504336 491668 504348
rect 483716 504308 491668 504336
rect 483716 504296 483722 504308
rect 491662 504296 491668 504308
rect 491720 504296 491726 504348
rect 512730 504296 512736 504348
rect 512788 504336 512794 504348
rect 519630 504336 519636 504348
rect 512788 504308 519636 504336
rect 512788 504296 512794 504308
rect 519630 504296 519636 504308
rect 519688 504296 519694 504348
rect 232682 504228 232688 504280
rect 232740 504268 232746 504280
rect 239766 504268 239772 504280
rect 232740 504240 239772 504268
rect 232740 504228 232746 504240
rect 239766 504228 239772 504240
rect 239824 504228 239830 504280
rect 316770 503752 316776 503804
rect 316828 503792 316834 503804
rect 323670 503792 323676 503804
rect 316828 503764 323676 503792
rect 316828 503752 316834 503764
rect 323670 503752 323676 503764
rect 323728 503752 323734 503804
rect 97902 503616 97908 503668
rect 97960 503656 97966 503668
rect 149054 503656 149060 503668
rect 97960 503628 149060 503656
rect 97960 503616 97966 503628
rect 149054 503616 149060 503628
rect 149112 503616 149118 503668
rect 182082 503616 182088 503668
rect 182140 503656 182146 503668
rect 233234 503656 233240 503668
rect 182140 503628 233240 503656
rect 182140 503616 182146 503628
rect 233234 503616 233240 503628
rect 233292 503616 233298 503668
rect 266262 503616 266268 503668
rect 266320 503656 266326 503668
rect 317414 503656 317420 503668
rect 266320 503628 317420 503656
rect 266320 503616 266326 503628
rect 317414 503616 317420 503628
rect 317472 503616 317478 503668
rect 378042 503616 378048 503668
rect 378100 503656 378106 503668
rect 429194 503656 429200 503668
rect 378100 503628 429200 503656
rect 378100 503616 378106 503628
rect 429194 503616 429200 503628
rect 429252 503616 429258 503668
rect 489822 503616 489828 503668
rect 489880 503656 489886 503668
rect 542354 503656 542360 503668
rect 489880 503628 542360 503656
rect 489880 503616 489886 503628
rect 542354 503616 542360 503628
rect 542412 503616 542418 503668
rect 427722 503548 427728 503600
rect 427780 503588 427786 503600
rect 428550 503588 428556 503600
rect 427780 503560 428556 503588
rect 427780 503548 427786 503560
rect 428550 503548 428556 503560
rect 428608 503548 428614 503600
rect 462222 503548 462228 503600
rect 462280 503588 462286 503600
rect 513374 503588 513380 503600
rect 462280 503560 513380 503588
rect 462280 503548 462286 503560
rect 513374 503548 513380 503560
rect 513432 503548 513438 503600
rect 35618 502256 35624 502308
rect 35676 502296 35682 502308
rect 36722 502296 36728 502308
rect 35676 502268 36728 502296
rect 35676 502256 35682 502268
rect 36722 502256 36728 502268
rect 36780 502256 36786 502308
rect 42886 500896 42892 500948
rect 42944 500936 42950 500948
rect 72050 500936 72056 500948
rect 42944 500908 45554 500936
rect 42944 500896 42950 500908
rect 15194 500828 15200 500880
rect 15252 500868 15258 500880
rect 43990 500868 43996 500880
rect 15252 500840 43996 500868
rect 15252 500828 15258 500840
rect 43990 500828 43996 500840
rect 44048 500828 44054 500880
rect 45526 500868 45554 500908
rect 64846 500908 72056 500936
rect 64846 500868 64874 500908
rect 72050 500896 72056 500908
rect 72108 500896 72114 500948
rect 99466 500896 99472 500948
rect 99524 500936 99530 500948
rect 99524 500908 103514 500936
rect 99524 500896 99530 500908
rect 45526 500840 64874 500868
rect 71866 500828 71872 500880
rect 71924 500868 71930 500880
rect 100018 500868 100024 500880
rect 71924 500840 100024 500868
rect 71924 500828 71930 500840
rect 100018 500828 100024 500840
rect 100076 500828 100082 500880
rect 103486 500868 103514 500908
rect 127066 500896 127072 500948
rect 127124 500936 127130 500948
rect 127124 500908 132494 500936
rect 127124 500896 127130 500908
rect 127986 500868 127992 500880
rect 103486 500840 127992 500868
rect 127986 500828 127992 500840
rect 128044 500828 128050 500880
rect 132466 500868 132494 500908
rect 183646 500896 183652 500948
rect 183704 500936 183710 500948
rect 183704 500908 190454 500936
rect 183704 500896 183710 500908
rect 156046 500868 156052 500880
rect 132466 500840 156052 500868
rect 156046 500828 156052 500840
rect 156104 500828 156110 500880
rect 165982 500828 165988 500880
rect 166040 500868 166046 500880
rect 177298 500868 177304 500880
rect 166040 500840 177304 500868
rect 166040 500828 166046 500840
rect 177298 500828 177304 500840
rect 177356 500828 177362 500880
rect 178678 500828 178684 500880
rect 178736 500868 178742 500880
rect 184014 500868 184020 500880
rect 178736 500840 184020 500868
rect 178736 500828 178742 500840
rect 184014 500828 184020 500840
rect 184072 500828 184078 500880
rect 190426 500868 190454 500908
rect 343358 500896 343364 500948
rect 343416 500936 343422 500948
rect 345658 500936 345664 500948
rect 343416 500908 345664 500936
rect 343416 500896 343422 500908
rect 345658 500896 345664 500908
rect 345716 500896 345722 500948
rect 374638 500896 374644 500948
rect 374696 500936 374702 500948
rect 379698 500936 379704 500948
rect 374696 500908 379704 500936
rect 374696 500896 374702 500908
rect 379698 500896 379704 500908
rect 379756 500896 379762 500948
rect 539318 500896 539324 500948
rect 539376 500936 539382 500948
rect 542998 500936 543004 500948
rect 539376 500908 543004 500936
rect 539376 500896 539382 500908
rect 542998 500896 543004 500908
rect 543056 500896 543062 500948
rect 211706 500868 211712 500880
rect 190426 500840 211712 500868
rect 211706 500828 211712 500840
rect 211764 500828 211770 500880
rect 222010 500828 222016 500880
rect 222068 500868 222074 500880
rect 232590 500868 232596 500880
rect 222068 500840 232596 500868
rect 222068 500828 222074 500840
rect 232590 500828 232596 500840
rect 232648 500828 232654 500880
rect 249702 500828 249708 500880
rect 249760 500868 249766 500880
rect 260098 500868 260104 500880
rect 249760 500840 260104 500868
rect 249760 500828 249766 500840
rect 260098 500828 260104 500840
rect 260156 500828 260162 500880
rect 261478 500828 261484 500880
rect 261536 500868 261542 500880
rect 567194 500868 567200 500880
rect 261536 500840 567200 500868
rect 261536 500828 261542 500840
rect 567194 500828 567200 500840
rect 567252 500828 567258 500880
rect 25682 500760 25688 500812
rect 25740 500800 25746 500812
rect 36998 500800 37004 500812
rect 25740 500772 37004 500800
rect 25740 500760 25746 500772
rect 36998 500760 37004 500772
rect 37056 500760 37062 500812
rect 53650 500760 53656 500812
rect 53708 500800 53714 500812
rect 69658 500800 69664 500812
rect 53708 500772 69664 500800
rect 53708 500760 53714 500772
rect 69658 500760 69664 500772
rect 69716 500760 69722 500812
rect 81986 500760 81992 500812
rect 82044 500800 82050 500812
rect 94498 500800 94504 500812
rect 82044 500772 94504 500800
rect 82044 500760 82050 500772
rect 94498 500760 94504 500772
rect 94556 500760 94562 500812
rect 109678 500760 109684 500812
rect 109736 500800 109742 500812
rect 120718 500800 120724 500812
rect 109736 500772 120724 500800
rect 109736 500760 109742 500772
rect 120718 500760 120724 500772
rect 120776 500760 120782 500812
rect 137646 500760 137652 500812
rect 137704 500800 137710 500812
rect 148318 500800 148324 500812
rect 137704 500772 148324 500800
rect 137704 500760 137710 500772
rect 148318 500760 148324 500772
rect 148376 500760 148382 500812
rect 193674 500760 193680 500812
rect 193732 500800 193738 500812
rect 204898 500800 204904 500812
rect 193732 500772 204904 500800
rect 193732 500760 193738 500772
rect 204898 500760 204904 500772
rect 204956 500760 204962 500812
rect 238846 500760 238852 500812
rect 238904 500800 238910 500812
rect 268010 500800 268016 500812
rect 238904 500772 268016 500800
rect 238904 500760 238910 500772
rect 268010 500760 268016 500772
rect 268068 500760 268074 500812
rect 277670 500760 277676 500812
rect 277728 500800 277734 500812
rect 289078 500800 289084 500812
rect 277728 500772 289084 500800
rect 277728 500760 277734 500772
rect 289078 500760 289084 500772
rect 289136 500760 289142 500812
rect 306006 500760 306012 500812
rect 306064 500800 306070 500812
rect 316678 500800 316684 500812
rect 306064 500772 316684 500800
rect 306064 500760 306070 500772
rect 316678 500760 316684 500772
rect 316736 500760 316742 500812
rect 323026 500760 323032 500812
rect 323084 500800 323090 500812
rect 352006 500800 352012 500812
rect 323084 500772 352012 500800
rect 323084 500760 323090 500772
rect 352006 500760 352012 500772
rect 352064 500760 352070 500812
rect 361666 500760 361672 500812
rect 361724 500800 361730 500812
rect 373258 500800 373264 500812
rect 361724 500772 373264 500800
rect 361724 500760 361730 500772
rect 373258 500760 373264 500772
rect 373316 500760 373322 500812
rect 379606 500760 379612 500812
rect 379664 500800 379670 500812
rect 408034 500800 408040 500812
rect 379664 500772 408040 500800
rect 379664 500760 379670 500772
rect 408034 500760 408040 500772
rect 408092 500760 408098 500812
rect 417694 500760 417700 500812
rect 417752 500800 417758 500812
rect 428458 500800 428464 500812
rect 417752 500772 428464 500800
rect 417752 500760 417758 500772
rect 428458 500760 428464 500772
rect 428516 500760 428522 500812
rect 434806 500760 434812 500812
rect 434864 500800 434870 500812
rect 463694 500800 463700 500812
rect 434864 500772 463700 500800
rect 434864 500760 434870 500772
rect 463694 500760 463700 500772
rect 463752 500760 463758 500812
rect 473998 500760 474004 500812
rect 474056 500800 474062 500812
rect 485038 500800 485044 500812
rect 474056 500772 485044 500800
rect 474056 500760 474062 500772
rect 485038 500760 485044 500772
rect 485096 500760 485102 500812
rect 501690 500760 501696 500812
rect 501748 500800 501754 500812
rect 512638 500800 512644 500812
rect 501748 500772 512644 500800
rect 501748 500760 501754 500772
rect 512638 500760 512644 500772
rect 512696 500760 512702 500812
rect 518986 500760 518992 500812
rect 519044 500800 519050 500812
rect 547874 500800 547880 500812
rect 519044 500772 547880 500800
rect 519044 500760 519050 500772
rect 547874 500760 547880 500772
rect 547932 500760 547938 500812
rect 333698 500692 333704 500744
rect 333756 500732 333762 500744
rect 344278 500732 344284 500744
rect 333756 500704 344284 500732
rect 333756 500692 333762 500704
rect 344278 500692 344284 500704
rect 344336 500692 344342 500744
rect 390002 500692 390008 500744
rect 390060 500732 390066 500744
rect 400858 500732 400864 500744
rect 390060 500704 400864 500732
rect 390060 500692 390066 500704
rect 400858 500692 400864 500704
rect 400916 500692 400922 500744
rect 445662 500692 445668 500744
rect 445720 500732 445726 500744
rect 456058 500732 456064 500744
rect 445720 500704 456064 500732
rect 445720 500692 445726 500704
rect 456058 500692 456064 500704
rect 456116 500692 456122 500744
rect 529658 500692 529664 500744
rect 529716 500732 529722 500744
rect 540238 500732 540244 500744
rect 529716 500704 540244 500732
rect 529716 500692 529722 500704
rect 540238 500692 540244 500704
rect 540296 500692 540302 500744
rect 36906 500624 36912 500676
rect 36964 500664 36970 500676
rect 557534 500664 557540 500676
rect 36964 500636 557540 500664
rect 36964 500624 36970 500636
rect 557534 500624 557540 500636
rect 557592 500624 557598 500676
rect 16022 497428 16028 497480
rect 16080 497468 16086 497480
rect 547874 497468 547880 497480
rect 16080 497440 547880 497468
rect 16080 497428 16086 497440
rect 547874 497428 547880 497440
rect 547932 497428 547938 497480
rect 25682 497088 25688 497140
rect 25740 497128 25746 497140
rect 261478 497128 261484 497140
rect 25740 497100 261484 497128
rect 25740 497088 25746 497100
rect 261478 497088 261484 497100
rect 261536 497088 261542 497140
rect 148410 497020 148416 497072
rect 148468 497060 148474 497072
rect 165706 497060 165712 497072
rect 148468 497032 165712 497060
rect 148468 497020 148474 497032
rect 165706 497020 165712 497032
rect 165764 497020 165770 497072
rect 175458 497020 175464 497072
rect 175516 497060 175522 497072
rect 193674 497060 193680 497072
rect 175516 497032 193680 497060
rect 175516 497020 175522 497032
rect 193674 497020 193680 497032
rect 193732 497020 193738 497072
rect 203518 497020 203524 497072
rect 203576 497060 203582 497072
rect 221366 497060 221372 497072
rect 203576 497032 221372 497060
rect 203576 497020 203582 497032
rect 221366 497020 221372 497032
rect 221424 497020 221430 497072
rect 408034 497020 408040 497072
rect 408092 497060 408098 497072
rect 428642 497060 428648 497072
rect 408092 497032 428648 497060
rect 408092 497020 408098 497032
rect 428642 497020 428648 497032
rect 428700 497020 428706 497072
rect 492030 497020 492036 497072
rect 492088 497060 492094 497072
rect 512730 497060 512736 497072
rect 492088 497032 512736 497060
rect 492088 497020 492094 497032
rect 512730 497020 512736 497032
rect 512788 497020 512794 497072
rect 36998 496952 37004 497004
rect 37056 496992 37062 497004
rect 53650 496992 53656 497004
rect 37056 496964 53656 496992
rect 37056 496952 37062 496964
rect 53650 496952 53656 496964
rect 53708 496952 53714 497004
rect 64322 496952 64328 497004
rect 64380 496992 64386 497004
rect 81434 496992 81440 497004
rect 64380 496964 81440 496992
rect 64380 496952 64386 496964
rect 81434 496952 81440 496964
rect 81492 496952 81498 497004
rect 91462 496952 91468 497004
rect 91520 496992 91526 497004
rect 109678 496992 109684 497004
rect 91520 496964 109684 496992
rect 91520 496952 91526 496964
rect 109678 496952 109684 496964
rect 109736 496952 109742 497004
rect 119430 496952 119436 497004
rect 119488 496992 119494 497004
rect 137646 496992 137652 497004
rect 119488 496964 137652 496992
rect 119488 496952 119494 496964
rect 137646 496952 137652 496964
rect 137704 496952 137710 497004
rect 156322 496952 156328 497004
rect 156380 496992 156386 497004
rect 178678 496992 178684 497004
rect 156380 496964 178684 496992
rect 156380 496952 156386 496964
rect 178678 496952 178684 496964
rect 178736 496952 178742 497004
rect 232498 496952 232504 497004
rect 232556 496992 232562 497004
rect 249702 496992 249708 497004
rect 232556 496964 249708 496992
rect 232556 496952 232562 496964
rect 249702 496952 249708 496964
rect 249760 496952 249766 497004
rect 260098 496952 260104 497004
rect 260156 496992 260162 497004
rect 277670 496992 277676 497004
rect 260156 496964 277676 496992
rect 260156 496952 260162 496964
rect 277670 496952 277676 496964
rect 277728 496952 277734 497004
rect 287514 496952 287520 497004
rect 287572 496992 287578 497004
rect 305362 496992 305368 497004
rect 287572 496964 305368 496992
rect 287572 496952 287578 496964
rect 305362 496952 305368 496964
rect 305420 496952 305426 497004
rect 315482 496952 315488 497004
rect 315540 496992 315546 497004
rect 333698 496992 333704 497004
rect 315540 496964 333704 496992
rect 315540 496952 315546 496964
rect 333698 496952 333704 496964
rect 333756 496952 333762 497004
rect 345658 496952 345664 497004
rect 345716 496992 345722 497004
rect 361666 496992 361672 497004
rect 345716 496964 361672 496992
rect 345716 496952 345722 496964
rect 361666 496952 361672 496964
rect 361724 496952 361730 497004
rect 371510 496952 371516 497004
rect 371568 496992 371574 497004
rect 389358 496992 389364 497004
rect 371568 496964 389364 496992
rect 371568 496952 371574 496964
rect 389358 496952 389364 496964
rect 389416 496952 389422 497004
rect 399478 496952 399484 497004
rect 399536 496992 399542 497004
rect 417694 496992 417700 497004
rect 399536 496964 417700 496992
rect 399536 496952 399542 496964
rect 417694 496952 417700 496964
rect 417752 496952 417758 497004
rect 456150 496952 456156 497004
rect 456208 496992 456214 497004
rect 473354 496992 473360 497004
rect 456208 496964 473360 496992
rect 456208 496952 456214 496964
rect 473354 496952 473360 496964
rect 473412 496952 473418 497004
rect 483474 496952 483480 497004
rect 483532 496992 483538 497004
rect 501690 496992 501696 497004
rect 483532 496964 501696 496992
rect 483532 496952 483538 496964
rect 501690 496952 501696 496964
rect 501748 496952 501754 497004
rect 36906 496884 36912 496936
rect 36964 496924 36970 496936
rect 63310 496924 63316 496936
rect 36964 496896 63316 496924
rect 36964 496884 36970 496896
rect 63310 496884 63316 496896
rect 63368 496884 63374 496936
rect 66898 496884 66904 496936
rect 66956 496924 66962 496936
rect 91094 496924 91100 496936
rect 66956 496896 91100 496924
rect 66956 496884 66962 496896
rect 91094 496884 91100 496896
rect 91152 496884 91158 496936
rect 94498 496884 94504 496936
rect 94556 496924 94562 496936
rect 119338 496924 119344 496936
rect 94556 496896 119344 496924
rect 94556 496884 94562 496896
rect 119338 496884 119344 496896
rect 119396 496884 119402 496936
rect 120718 496884 120724 496936
rect 120776 496924 120782 496936
rect 147306 496924 147312 496936
rect 120776 496896 147312 496924
rect 120776 496884 120782 496896
rect 147306 496884 147312 496896
rect 147364 496884 147370 496936
rect 148318 496884 148324 496936
rect 148376 496924 148382 496936
rect 175366 496924 175372 496936
rect 148376 496896 175372 496924
rect 148376 496884 148382 496896
rect 175366 496884 175372 496896
rect 175424 496884 175430 496936
rect 177298 496884 177304 496936
rect 177356 496924 177362 496936
rect 203334 496924 203340 496936
rect 177356 496896 203340 496924
rect 177356 496884 177362 496896
rect 203334 496884 203340 496896
rect 203392 496884 203398 496936
rect 204898 496884 204904 496936
rect 204956 496924 204962 496936
rect 231026 496924 231032 496936
rect 204956 496896 231032 496924
rect 204956 496884 204962 496896
rect 231026 496884 231032 496896
rect 231084 496884 231090 496936
rect 232590 496884 232596 496936
rect 232648 496924 232654 496936
rect 259362 496924 259368 496936
rect 232648 496896 259368 496924
rect 232648 496884 232654 496896
rect 259362 496884 259368 496896
rect 259420 496884 259426 496936
rect 268010 496884 268016 496936
rect 268068 496924 268074 496936
rect 287698 496924 287704 496936
rect 268068 496896 287704 496924
rect 268068 496884 268074 496896
rect 287698 496884 287704 496896
rect 287756 496884 287762 496936
rect 296346 496884 296352 496936
rect 296404 496924 296410 496936
rect 316770 496924 316776 496936
rect 296404 496896 316776 496924
rect 296404 496884 296410 496896
rect 316770 496884 316776 496896
rect 316828 496884 316834 496936
rect 352006 496884 352012 496936
rect 352064 496924 352070 496936
rect 374638 496924 374644 496936
rect 352064 496896 374644 496924
rect 352064 496884 352070 496896
rect 374638 496884 374644 496896
rect 374696 496884 374702 496936
rect 428550 496884 428556 496936
rect 428608 496924 428614 496936
rect 445662 496924 445668 496936
rect 428608 496896 445668 496924
rect 428608 496884 428614 496896
rect 445662 496884 445668 496896
rect 445720 496884 445726 496936
rect 464338 496884 464344 496936
rect 464396 496924 464402 496936
rect 483658 496924 483664 496936
rect 464396 496896 483664 496924
rect 464396 496884 464402 496896
rect 483658 496884 483664 496896
rect 483716 496884 483722 496936
rect 511442 496884 511448 496936
rect 511500 496924 511506 496936
rect 529658 496924 529664 496936
rect 511500 496896 529664 496924
rect 511500 496884 511506 496896
rect 529658 496884 529664 496896
rect 529716 496884 529722 496936
rect 542998 496884 543004 496936
rect 543056 496924 543062 496936
rect 557534 496924 557540 496936
rect 543056 496896 557540 496924
rect 543056 496884 543062 496896
rect 557534 496884 557540 496896
rect 557592 496884 557598 496936
rect 212350 496816 212356 496868
rect 212408 496856 212414 496868
rect 232682 496856 232688 496868
rect 212408 496828 232688 496856
rect 212408 496816 212414 496828
rect 232682 496816 232688 496828
rect 232740 496816 232746 496868
rect 260190 496816 260196 496868
rect 260248 496856 260254 496868
rect 287330 496856 287336 496868
rect 260248 496828 287336 496856
rect 260248 496816 260254 496828
rect 287330 496816 287336 496828
rect 287388 496816 287394 496868
rect 289078 496816 289084 496868
rect 289136 496856 289142 496868
rect 315022 496856 315028 496868
rect 289136 496828 315028 496856
rect 289136 496816 289142 496828
rect 315022 496816 315028 496828
rect 315080 496816 315086 496868
rect 316678 496816 316684 496868
rect 316736 496856 316742 496868
rect 343358 496856 343364 496868
rect 316736 496828 343364 496856
rect 316736 496816 316742 496828
rect 343358 496816 343364 496828
rect 343416 496816 343422 496868
rect 344278 496816 344284 496868
rect 344336 496856 344342 496868
rect 371326 496856 371332 496868
rect 344336 496828 371332 496856
rect 344336 496816 344342 496828
rect 371326 496816 371332 496828
rect 371384 496816 371390 496868
rect 373258 496816 373264 496868
rect 373316 496856 373322 496868
rect 399018 496856 399024 496868
rect 373316 496828 399024 496856
rect 373316 496816 373322 496828
rect 399018 496816 399024 496828
rect 399076 496816 399082 496868
rect 400858 496816 400864 496868
rect 400916 496856 400922 496868
rect 427354 496856 427360 496868
rect 400916 496828 427360 496856
rect 400916 496816 400922 496828
rect 427354 496816 427360 496828
rect 427412 496816 427418 496868
rect 428458 496816 428464 496868
rect 428516 496856 428522 496868
rect 455322 496856 455328 496868
rect 428516 496828 455328 496856
rect 428516 496816 428522 496828
rect 455322 496816 455328 496828
rect 455380 496816 455386 496868
rect 456058 496816 456064 496868
rect 456116 496856 456122 496868
rect 483014 496856 483020 496868
rect 456116 496828 483020 496856
rect 456116 496816 456122 496828
rect 483014 496816 483020 496828
rect 483072 496816 483078 496868
rect 485038 496816 485044 496868
rect 485096 496856 485102 496868
rect 511350 496856 511356 496868
rect 485096 496828 511356 496856
rect 485096 496816 485102 496828
rect 511350 496816 511356 496828
rect 511408 496816 511414 496868
rect 512638 496816 512644 496868
rect 512696 496856 512702 496868
rect 539318 496856 539324 496868
rect 512696 496828 539324 496856
rect 512696 496816 512702 496828
rect 539318 496816 539324 496828
rect 539376 496816 539382 496868
rect 540238 496816 540244 496868
rect 540296 496856 540302 496868
rect 567194 496856 567200 496868
rect 540296 496828 567200 496856
rect 540296 496816 540302 496828
rect 567194 496816 567200 496828
rect 567252 496816 567258 496868
rect 37918 494708 37924 494760
rect 37976 494748 37982 494760
rect 545758 494748 545764 494760
rect 37976 494720 545764 494748
rect 37976 494708 37982 494720
rect 545758 494708 545764 494720
rect 545816 494708 545822 494760
rect 35618 494028 35624 494080
rect 35676 494068 35682 494080
rect 36722 494068 36728 494080
rect 35676 494040 36728 494068
rect 35676 494028 35682 494040
rect 36722 494028 36728 494040
rect 36780 494028 36786 494080
rect 63586 477640 63592 477692
rect 63644 477680 63650 477692
rect 64322 477680 64328 477692
rect 63644 477652 64328 477680
rect 63644 477640 63650 477652
rect 64322 477640 64328 477652
rect 64380 477640 64386 477692
rect 147674 477640 147680 477692
rect 147732 477680 147738 477692
rect 148410 477680 148416 477692
rect 147732 477652 148416 477680
rect 147732 477640 147738 477652
rect 148410 477640 148416 477652
rect 148468 477640 148474 477692
rect 455690 477640 455696 477692
rect 455748 477680 455754 477692
rect 456150 477680 456156 477692
rect 455748 477652 456156 477680
rect 455748 477640 455754 477652
rect 456150 477640 456156 477652
rect 456208 477640 456214 477692
rect 512730 476960 512736 477012
rect 512788 477000 512794 477012
rect 519630 477000 519636 477012
rect 512788 476972 519636 477000
rect 512788 476960 512794 476972
rect 519630 476960 519636 476972
rect 519688 476960 519694 477012
rect 428642 476756 428648 476808
rect 428700 476796 428706 476808
rect 435726 476796 435732 476808
rect 428700 476768 435732 476796
rect 428700 476756 428706 476768
rect 435726 476756 435732 476768
rect 435784 476756 435790 476808
rect 232682 476552 232688 476604
rect 232740 476592 232746 476604
rect 239766 476592 239772 476604
rect 232740 476564 239772 476592
rect 232740 476552 232746 476564
rect 239766 476552 239772 476564
rect 239824 476552 239830 476604
rect 287698 476416 287704 476468
rect 287756 476456 287762 476468
rect 295702 476456 295708 476468
rect 287756 476428 295708 476456
rect 287756 476416 287762 476428
rect 295702 476416 295708 476428
rect 295760 476416 295766 476468
rect 316770 476416 316776 476468
rect 316828 476456 316834 476468
rect 323670 476456 323676 476468
rect 316828 476428 323676 476456
rect 316828 476416 316834 476428
rect 323670 476416 323676 476428
rect 323728 476416 323734 476468
rect 483658 476280 483664 476332
rect 483716 476320 483722 476332
rect 491662 476320 491668 476332
rect 483716 476292 491668 476320
rect 483716 476280 483722 476292
rect 491662 476280 491668 476292
rect 491720 476280 491726 476332
rect 13722 476008 13728 476060
rect 13780 476048 13786 476060
rect 66254 476048 66260 476060
rect 13780 476020 66260 476048
rect 13780 476008 13786 476020
rect 66254 476008 66260 476020
rect 66312 476008 66318 476060
rect 70302 476008 70308 476060
rect 70360 476048 70366 476060
rect 121454 476048 121460 476060
rect 70360 476020 121460 476048
rect 70360 476008 70366 476020
rect 121454 476008 121460 476020
rect 121512 476008 121518 476060
rect 126882 476008 126888 476060
rect 126940 476048 126946 476060
rect 178034 476048 178040 476060
rect 126940 476020 178040 476048
rect 126940 476008 126946 476020
rect 178034 476008 178040 476020
rect 178092 476008 178098 476060
rect 209682 476008 209688 476060
rect 209740 476048 209746 476060
rect 262214 476048 262220 476060
rect 209740 476020 262220 476048
rect 209740 476008 209746 476020
rect 262214 476008 262220 476020
rect 262272 476008 262278 476060
rect 266262 476008 266268 476060
rect 266320 476048 266326 476060
rect 317414 476048 317420 476060
rect 266320 476020 317420 476048
rect 266320 476008 266326 476020
rect 317414 476008 317420 476020
rect 317472 476008 317478 476060
rect 322842 476008 322848 476060
rect 322900 476048 322906 476060
rect 373994 476048 374000 476060
rect 322900 476020 374000 476048
rect 322900 476008 322906 476020
rect 373994 476008 374000 476020
rect 374052 476008 374058 476060
rect 405642 476008 405648 476060
rect 405700 476048 405706 476060
rect 458174 476048 458180 476060
rect 405700 476020 458180 476048
rect 405700 476008 405706 476020
rect 458174 476008 458180 476020
rect 458232 476008 458238 476060
rect 489822 476008 489828 476060
rect 489880 476048 489886 476060
rect 542354 476048 542360 476060
rect 489880 476020 542360 476048
rect 489880 476008 489886 476020
rect 542354 476008 542360 476020
rect 542412 476008 542418 476060
rect 35618 475940 35624 475992
rect 35676 475980 35682 475992
rect 36998 475980 37004 475992
rect 35676 475952 37004 475980
rect 35676 475940 35682 475952
rect 36998 475940 37004 475952
rect 37056 475940 37062 475992
rect 42702 475940 42708 475992
rect 42760 475980 42766 475992
rect 93854 475980 93860 475992
rect 42760 475952 93860 475980
rect 42760 475940 42766 475952
rect 93854 475940 93860 475952
rect 93912 475940 93918 475992
rect 97902 475940 97908 475992
rect 97960 475980 97966 475992
rect 149054 475980 149060 475992
rect 97960 475952 149060 475980
rect 97960 475940 97966 475952
rect 149054 475940 149060 475952
rect 149112 475940 149118 475992
rect 154482 475940 154488 475992
rect 154540 475980 154546 475992
rect 205634 475980 205640 475992
rect 154540 475952 205640 475980
rect 154540 475940 154546 475952
rect 205634 475940 205640 475952
rect 205692 475940 205698 475992
rect 238662 475940 238668 475992
rect 238720 475980 238726 475992
rect 289814 475980 289820 475992
rect 238720 475952 289820 475980
rect 238720 475940 238726 475952
rect 289814 475940 289820 475952
rect 289872 475940 289878 475992
rect 293862 475940 293868 475992
rect 293920 475980 293926 475992
rect 345014 475980 345020 475992
rect 293920 475952 345020 475980
rect 293920 475940 293926 475952
rect 345014 475940 345020 475952
rect 345072 475940 345078 475992
rect 350442 475940 350448 475992
rect 350500 475980 350506 475992
rect 401594 475980 401600 475992
rect 350500 475952 401600 475980
rect 350500 475940 350506 475952
rect 401594 475940 401600 475952
rect 401652 475940 401658 475992
rect 427722 475940 427728 475992
rect 427780 475980 427786 475992
rect 428550 475980 428556 475992
rect 427780 475952 428556 475980
rect 427780 475940 427786 475952
rect 428550 475940 428556 475952
rect 428608 475940 428614 475992
rect 434622 475940 434628 475992
rect 434680 475980 434686 475992
rect 485774 475980 485780 475992
rect 434680 475952 485780 475980
rect 434680 475940 434686 475952
rect 485774 475940 485780 475952
rect 485832 475940 485838 475992
rect 518802 475940 518808 475992
rect 518860 475980 518866 475992
rect 569954 475980 569960 475992
rect 518860 475952 569960 475980
rect 518860 475940 518866 475952
rect 569954 475940 569960 475952
rect 570012 475940 570018 475992
rect 182082 475872 182088 475924
rect 182140 475912 182146 475924
rect 233234 475912 233240 475924
rect 182140 475884 233240 475912
rect 182140 475872 182146 475884
rect 233234 475872 233240 475884
rect 233292 475872 233298 475924
rect 343542 475872 343548 475924
rect 343600 475912 343606 475924
rect 345658 475912 345664 475924
rect 343600 475884 345664 475912
rect 343600 475872 343606 475884
rect 345658 475872 345664 475884
rect 345716 475872 345722 475924
rect 378042 475872 378048 475924
rect 378100 475912 378106 475924
rect 429194 475912 429200 475924
rect 378100 475884 429200 475912
rect 378100 475872 378106 475884
rect 429194 475872 429200 475884
rect 429252 475872 429258 475924
rect 462222 475872 462228 475924
rect 462280 475912 462286 475924
rect 513374 475912 513380 475924
rect 462280 475884 513380 475912
rect 462280 475872 462286 475884
rect 513374 475872 513380 475884
rect 513432 475872 513438 475924
rect 539502 475872 539508 475924
rect 539560 475912 539566 475924
rect 542998 475912 543004 475924
rect 539560 475884 543004 475912
rect 539560 475872 539566 475884
rect 542998 475872 543004 475884
rect 543056 475872 543062 475924
rect 178678 473288 178684 473340
rect 178736 473328 178742 473340
rect 184014 473328 184020 473340
rect 178736 473300 184020 473328
rect 178736 473288 178742 473300
rect 184014 473288 184020 473300
rect 184072 473288 184078 473340
rect 374638 473288 374644 473340
rect 374696 473328 374702 473340
rect 379698 473328 379704 473340
rect 374696 473300 379704 473328
rect 374696 473288 374702 473300
rect 379698 473288 379704 473300
rect 379756 473288 379762 473340
rect 15194 473220 15200 473272
rect 15252 473260 15258 473272
rect 43990 473260 43996 473272
rect 15252 473232 43996 473260
rect 15252 473220 15258 473232
rect 43990 473220 43996 473232
rect 44048 473220 44054 473272
rect 71038 473220 71044 473272
rect 71096 473260 71102 473272
rect 567194 473260 567200 473272
rect 71096 473232 567200 473260
rect 71096 473220 71102 473232
rect 567194 473220 567200 473232
rect 567252 473220 567258 473272
rect 25682 473152 25688 473204
rect 25740 473192 25746 473204
rect 36906 473192 36912 473204
rect 25740 473164 36912 473192
rect 25740 473152 25746 473164
rect 36906 473152 36912 473164
rect 36964 473152 36970 473204
rect 53650 473152 53656 473204
rect 53708 473192 53714 473204
rect 66898 473192 66904 473204
rect 53708 473164 66904 473192
rect 53708 473152 53714 473164
rect 66898 473152 66904 473164
rect 66956 473152 66962 473204
rect 71866 473152 71872 473204
rect 71924 473192 71930 473204
rect 100018 473192 100024 473204
rect 71924 473164 100024 473192
rect 71924 473152 71930 473164
rect 100018 473152 100024 473164
rect 100076 473152 100082 473204
rect 127986 473192 127992 473204
rect 103486 473164 127992 473192
rect 42886 473084 42892 473136
rect 42944 473124 42950 473136
rect 72050 473124 72056 473136
rect 42944 473096 72056 473124
rect 42944 473084 42950 473096
rect 72050 473084 72056 473096
rect 72108 473084 72114 473136
rect 81986 473084 81992 473136
rect 82044 473124 82050 473136
rect 94498 473124 94504 473136
rect 82044 473096 94504 473124
rect 82044 473084 82050 473096
rect 94498 473084 94504 473096
rect 94556 473084 94562 473136
rect 99466 473084 99472 473136
rect 99524 473124 99530 473136
rect 103486 473124 103514 473164
rect 127986 473152 127992 473164
rect 128044 473152 128050 473204
rect 156046 473192 156052 473204
rect 132466 473164 156052 473192
rect 99524 473096 103514 473124
rect 99524 473084 99530 473096
rect 109678 473084 109684 473136
rect 109736 473124 109742 473136
rect 120718 473124 120724 473136
rect 109736 473096 120724 473124
rect 109736 473084 109742 473096
rect 120718 473084 120724 473096
rect 120776 473084 120782 473136
rect 127066 473084 127072 473136
rect 127124 473124 127130 473136
rect 132466 473124 132494 473164
rect 156046 473152 156052 473164
rect 156104 473152 156110 473204
rect 165982 473152 165988 473204
rect 166040 473192 166046 473204
rect 177298 473192 177304 473204
rect 166040 473164 177304 473192
rect 166040 473152 166046 473164
rect 177298 473152 177304 473164
rect 177356 473152 177362 473204
rect 183646 473152 183652 473204
rect 183704 473192 183710 473204
rect 211706 473192 211712 473204
rect 183704 473164 211712 473192
rect 183704 473152 183710 473164
rect 211706 473152 211712 473164
rect 211764 473152 211770 473204
rect 222010 473152 222016 473204
rect 222068 473192 222074 473204
rect 232590 473192 232596 473204
rect 222068 473164 232596 473192
rect 222068 473152 222074 473164
rect 232590 473152 232596 473164
rect 232648 473152 232654 473204
rect 238846 473152 238852 473204
rect 238904 473192 238910 473204
rect 268010 473192 268016 473204
rect 238904 473164 268016 473192
rect 238904 473152 238910 473164
rect 268010 473152 268016 473164
rect 268068 473152 268074 473204
rect 277670 473152 277676 473204
rect 277728 473192 277734 473204
rect 289078 473192 289084 473204
rect 277728 473164 289084 473192
rect 277728 473152 277734 473164
rect 289078 473152 289084 473164
rect 289136 473152 289142 473204
rect 306006 473152 306012 473204
rect 306064 473192 306070 473204
rect 316678 473192 316684 473204
rect 306064 473164 316684 473192
rect 306064 473152 306070 473164
rect 316678 473152 316684 473164
rect 316736 473152 316742 473204
rect 323026 473152 323032 473204
rect 323084 473192 323090 473204
rect 352006 473192 352012 473204
rect 323084 473164 352012 473192
rect 323084 473152 323090 473164
rect 352006 473152 352012 473164
rect 352064 473152 352070 473204
rect 361666 473152 361672 473204
rect 361724 473192 361730 473204
rect 373258 473192 373264 473204
rect 361724 473164 373264 473192
rect 361724 473152 361730 473164
rect 373258 473152 373264 473164
rect 373316 473152 373322 473204
rect 379606 473152 379612 473204
rect 379664 473192 379670 473204
rect 408034 473192 408040 473204
rect 379664 473164 408040 473192
rect 379664 473152 379670 473164
rect 408034 473152 408040 473164
rect 408092 473152 408098 473204
rect 417694 473152 417700 473204
rect 417752 473192 417758 473204
rect 428458 473192 428464 473204
rect 417752 473164 428464 473192
rect 417752 473152 417758 473164
rect 428458 473152 428464 473164
rect 428516 473152 428522 473204
rect 434806 473152 434812 473204
rect 434864 473192 434870 473204
rect 463694 473192 463700 473204
rect 434864 473164 463700 473192
rect 434864 473152 434870 473164
rect 463694 473152 463700 473164
rect 463752 473152 463758 473204
rect 473998 473152 474004 473204
rect 474056 473192 474062 473204
rect 485038 473192 485044 473204
rect 474056 473164 485044 473192
rect 474056 473152 474062 473164
rect 485038 473152 485044 473164
rect 485096 473152 485102 473204
rect 501690 473152 501696 473204
rect 501748 473192 501754 473204
rect 512638 473192 512644 473204
rect 501748 473164 512644 473192
rect 501748 473152 501754 473164
rect 512638 473152 512644 473164
rect 512696 473152 512702 473204
rect 518986 473152 518992 473204
rect 519044 473192 519050 473204
rect 547874 473192 547880 473204
rect 519044 473164 547880 473192
rect 519044 473152 519050 473164
rect 547874 473152 547880 473164
rect 547932 473152 547938 473204
rect 127124 473096 132494 473124
rect 127124 473084 127130 473096
rect 137646 473084 137652 473136
rect 137704 473124 137710 473136
rect 148318 473124 148324 473136
rect 137704 473096 148324 473124
rect 137704 473084 137710 473096
rect 148318 473084 148324 473096
rect 148376 473084 148382 473136
rect 193674 473084 193680 473136
rect 193732 473124 193738 473136
rect 204898 473124 204904 473136
rect 193732 473096 204904 473124
rect 193732 473084 193738 473096
rect 204898 473084 204904 473096
rect 204956 473084 204962 473136
rect 249702 473084 249708 473136
rect 249760 473124 249766 473136
rect 260190 473124 260196 473136
rect 249760 473096 260196 473124
rect 249760 473084 249766 473096
rect 260190 473084 260196 473096
rect 260248 473084 260254 473136
rect 333698 473084 333704 473136
rect 333756 473124 333762 473136
rect 344278 473124 344284 473136
rect 333756 473096 344284 473124
rect 333756 473084 333762 473096
rect 344278 473084 344284 473096
rect 344336 473084 344342 473136
rect 390002 473084 390008 473136
rect 390060 473124 390066 473136
rect 400858 473124 400864 473136
rect 390060 473096 400864 473124
rect 390060 473084 390066 473096
rect 400858 473084 400864 473096
rect 400916 473084 400922 473136
rect 445662 473084 445668 473136
rect 445720 473124 445726 473136
rect 456058 473124 456064 473136
rect 445720 473096 456064 473124
rect 445720 473084 445726 473096
rect 456058 473084 456064 473096
rect 456116 473084 456122 473136
rect 529658 473084 529664 473136
rect 529716 473124 529722 473136
rect 540238 473124 540244 473136
rect 529716 473096 540244 473124
rect 529716 473084 529722 473096
rect 540238 473084 540244 473096
rect 540296 473084 540302 473136
rect 36814 473016 36820 473068
rect 36872 473056 36878 473068
rect 557534 473056 557540 473068
rect 36872 473028 557540 473056
rect 36872 473016 36878 473028
rect 557534 473016 557540 473028
rect 557592 473016 557598 473068
rect 15286 469820 15292 469872
rect 15344 469860 15350 469872
rect 547874 469860 547880 469872
rect 15344 469832 547880 469860
rect 15344 469820 15350 469832
rect 547874 469820 547880 469832
rect 547932 469820 547938 469872
rect 25682 469412 25688 469464
rect 25740 469452 25746 469464
rect 71038 469452 71044 469464
rect 25740 469424 71044 469452
rect 25740 469412 25746 469424
rect 71038 469412 71044 469424
rect 71096 469412 71102 469464
rect 296346 469412 296352 469464
rect 296404 469452 296410 469464
rect 316770 469452 316776 469464
rect 296404 469424 316776 469452
rect 296404 469412 296410 469424
rect 316770 469412 316776 469424
rect 316828 469412 316834 469464
rect 408034 469412 408040 469464
rect 408092 469452 408098 469464
rect 428642 469452 428648 469464
rect 408092 469424 428648 469452
rect 408092 469412 408098 469424
rect 428642 469412 428648 469424
rect 428700 469412 428706 469464
rect 36998 469344 37004 469396
rect 37056 469384 37062 469396
rect 53650 469384 53656 469396
rect 37056 469356 53656 469384
rect 37056 469344 37062 469356
rect 53650 469344 53656 469356
rect 53708 469344 53714 469396
rect 148410 469344 148416 469396
rect 148468 469384 148474 469396
rect 165706 469384 165712 469396
rect 148468 469356 165712 469384
rect 148468 469344 148474 469356
rect 165706 469344 165712 469356
rect 165764 469344 165770 469396
rect 175458 469344 175464 469396
rect 175516 469384 175522 469396
rect 193674 469384 193680 469396
rect 175516 469356 193680 469384
rect 175516 469344 175522 469356
rect 193674 469344 193680 469356
rect 193732 469344 193738 469396
rect 203518 469344 203524 469396
rect 203576 469384 203582 469396
rect 221366 469384 221372 469396
rect 203576 469356 221372 469384
rect 203576 469344 203582 469356
rect 221366 469344 221372 469356
rect 221424 469344 221430 469396
rect 232498 469344 232504 469396
rect 232556 469384 232562 469396
rect 249702 469384 249708 469396
rect 232556 469356 249708 469384
rect 232556 469344 232562 469356
rect 249702 469344 249708 469356
rect 249760 469344 249766 469396
rect 260098 469344 260104 469396
rect 260156 469384 260162 469396
rect 277670 469384 277676 469396
rect 260156 469356 277676 469384
rect 260156 469344 260162 469356
rect 277670 469344 277676 469356
rect 277728 469344 277734 469396
rect 287514 469344 287520 469396
rect 287572 469384 287578 469396
rect 305362 469384 305368 469396
rect 287572 469356 305368 469384
rect 287572 469344 287578 469356
rect 305362 469344 305368 469356
rect 305420 469344 305426 469396
rect 345658 469344 345664 469396
rect 345716 469384 345722 469396
rect 361666 469384 361672 469396
rect 345716 469356 361672 469384
rect 345716 469344 345722 469356
rect 361666 469344 361672 469356
rect 361724 469344 361730 469396
rect 371510 469344 371516 469396
rect 371568 469384 371574 469396
rect 389358 469384 389364 469396
rect 371568 469356 389364 469384
rect 371568 469344 371574 469356
rect 389358 469344 389364 469356
rect 389416 469344 389422 469396
rect 399478 469344 399484 469396
rect 399536 469384 399542 469396
rect 417694 469384 417700 469396
rect 399536 469356 417700 469384
rect 399536 469344 399542 469356
rect 417694 469344 417700 469356
rect 417752 469344 417758 469396
rect 456150 469344 456156 469396
rect 456208 469384 456214 469396
rect 473354 469384 473360 469396
rect 456208 469356 473360 469384
rect 456208 469344 456214 469356
rect 473354 469344 473360 469356
rect 473412 469344 473418 469396
rect 483474 469344 483480 469396
rect 483532 469384 483538 469396
rect 501690 469384 501696 469396
rect 483532 469356 501696 469384
rect 483532 469344 483538 469356
rect 501690 469344 501696 469356
rect 501748 469344 501754 469396
rect 511442 469344 511448 469396
rect 511500 469384 511506 469396
rect 529658 469384 529664 469396
rect 511500 469356 529664 469384
rect 511500 469344 511506 469356
rect 529658 469344 529664 469356
rect 529716 469344 529722 469396
rect 36906 469276 36912 469328
rect 36964 469316 36970 469328
rect 63310 469316 63316 469328
rect 36964 469288 63316 469316
rect 36964 469276 36970 469288
rect 63310 469276 63316 469288
rect 63368 469276 63374 469328
rect 64322 469276 64328 469328
rect 64380 469316 64386 469328
rect 81434 469316 81440 469328
rect 64380 469288 81440 469316
rect 64380 469276 64386 469288
rect 81434 469276 81440 469288
rect 81492 469276 81498 469328
rect 91462 469276 91468 469328
rect 91520 469316 91526 469328
rect 109678 469316 109684 469328
rect 91520 469288 109684 469316
rect 91520 469276 91526 469288
rect 109678 469276 109684 469288
rect 109736 469276 109742 469328
rect 119430 469276 119436 469328
rect 119488 469316 119494 469328
rect 137646 469316 137652 469328
rect 119488 469288 137652 469316
rect 119488 469276 119494 469288
rect 137646 469276 137652 469288
rect 137704 469276 137710 469328
rect 156322 469276 156328 469328
rect 156380 469316 156386 469328
rect 178678 469316 178684 469328
rect 156380 469288 178684 469316
rect 156380 469276 156386 469288
rect 178678 469276 178684 469288
rect 178736 469276 178742 469328
rect 212350 469276 212356 469328
rect 212408 469316 212414 469328
rect 232682 469316 232688 469328
rect 212408 469288 232688 469316
rect 212408 469276 212414 469288
rect 232682 469276 232688 469288
rect 232740 469276 232746 469328
rect 268010 469276 268016 469328
rect 268068 469316 268074 469328
rect 287698 469316 287704 469328
rect 268068 469288 287704 469316
rect 268068 469276 268074 469288
rect 287698 469276 287704 469288
rect 287756 469276 287762 469328
rect 315482 469276 315488 469328
rect 315540 469316 315546 469328
rect 333698 469316 333704 469328
rect 315540 469288 333704 469316
rect 315540 469276 315546 469288
rect 333698 469276 333704 469288
rect 333756 469276 333762 469328
rect 352006 469276 352012 469328
rect 352064 469316 352070 469328
rect 374638 469316 374644 469328
rect 352064 469288 374644 469316
rect 352064 469276 352070 469288
rect 374638 469276 374644 469288
rect 374696 469276 374702 469328
rect 428458 469276 428464 469328
rect 428516 469316 428522 469328
rect 445662 469316 445668 469328
rect 428516 469288 445668 469316
rect 428516 469276 428522 469288
rect 445662 469276 445668 469288
rect 445720 469276 445726 469328
rect 464338 469276 464344 469328
rect 464396 469316 464402 469328
rect 483658 469316 483664 469328
rect 464396 469288 483664 469316
rect 464396 469276 464402 469288
rect 483658 469276 483664 469288
rect 483716 469276 483722 469328
rect 492030 469276 492036 469328
rect 492088 469316 492094 469328
rect 512730 469316 512736 469328
rect 492088 469288 512736 469316
rect 492088 469276 492094 469288
rect 512730 469276 512736 469288
rect 512788 469276 512794 469328
rect 542998 469276 543004 469328
rect 543056 469316 543062 469328
rect 557534 469316 557540 469328
rect 543056 469288 557540 469316
rect 543056 469276 543062 469288
rect 557534 469276 557540 469288
rect 557592 469276 557598 469328
rect 69658 469208 69664 469260
rect 69716 469248 69722 469260
rect 91094 469248 91100 469260
rect 69716 469220 91100 469248
rect 69716 469208 69722 469220
rect 91094 469208 91100 469220
rect 91152 469208 91158 469260
rect 94498 469208 94504 469260
rect 94556 469248 94562 469260
rect 119338 469248 119344 469260
rect 94556 469220 119344 469248
rect 94556 469208 94562 469220
rect 119338 469208 119344 469220
rect 119396 469208 119402 469260
rect 120718 469208 120724 469260
rect 120776 469248 120782 469260
rect 147306 469248 147312 469260
rect 120776 469220 147312 469248
rect 120776 469208 120782 469220
rect 147306 469208 147312 469220
rect 147364 469208 147370 469260
rect 148318 469208 148324 469260
rect 148376 469248 148382 469260
rect 175366 469248 175372 469260
rect 148376 469220 175372 469248
rect 148376 469208 148382 469220
rect 175366 469208 175372 469220
rect 175424 469208 175430 469260
rect 177298 469208 177304 469260
rect 177356 469248 177362 469260
rect 203334 469248 203340 469260
rect 177356 469220 203340 469248
rect 177356 469208 177362 469220
rect 203334 469208 203340 469220
rect 203392 469208 203398 469260
rect 204898 469208 204904 469260
rect 204956 469248 204962 469260
rect 231026 469248 231032 469260
rect 204956 469220 231032 469248
rect 204956 469208 204962 469220
rect 231026 469208 231032 469220
rect 231084 469208 231090 469260
rect 232590 469208 232596 469260
rect 232648 469248 232654 469260
rect 259362 469248 259368 469260
rect 232648 469220 259368 469248
rect 232648 469208 232654 469220
rect 259362 469208 259368 469220
rect 259420 469208 259426 469260
rect 260190 469208 260196 469260
rect 260248 469248 260254 469260
rect 287330 469248 287336 469260
rect 260248 469220 287336 469248
rect 260248 469208 260254 469220
rect 287330 469208 287336 469220
rect 287388 469208 287394 469260
rect 289078 469208 289084 469260
rect 289136 469248 289142 469260
rect 315022 469248 315028 469260
rect 289136 469220 315028 469248
rect 289136 469208 289142 469220
rect 315022 469208 315028 469220
rect 315080 469208 315086 469260
rect 316678 469208 316684 469260
rect 316736 469248 316742 469260
rect 343358 469248 343364 469260
rect 316736 469220 343364 469248
rect 316736 469208 316742 469220
rect 343358 469208 343364 469220
rect 343416 469208 343422 469260
rect 344278 469208 344284 469260
rect 344336 469248 344342 469260
rect 371326 469248 371332 469260
rect 344336 469220 371332 469248
rect 344336 469208 344342 469220
rect 371326 469208 371332 469220
rect 371384 469208 371390 469260
rect 373258 469208 373264 469260
rect 373316 469248 373322 469260
rect 399018 469248 399024 469260
rect 373316 469220 399024 469248
rect 373316 469208 373322 469220
rect 399018 469208 399024 469220
rect 399076 469208 399082 469260
rect 400858 469208 400864 469260
rect 400916 469248 400922 469260
rect 427354 469248 427360 469260
rect 400916 469220 427360 469248
rect 400916 469208 400922 469220
rect 427354 469208 427360 469220
rect 427412 469208 427418 469260
rect 428550 469208 428556 469260
rect 428608 469248 428614 469260
rect 455322 469248 455328 469260
rect 428608 469220 455328 469248
rect 428608 469208 428614 469220
rect 455322 469208 455328 469220
rect 455380 469208 455386 469260
rect 456058 469208 456064 469260
rect 456116 469248 456122 469260
rect 483014 469248 483020 469260
rect 456116 469220 483020 469248
rect 456116 469208 456122 469220
rect 483014 469208 483020 469220
rect 483072 469208 483078 469260
rect 485038 469208 485044 469260
rect 485096 469248 485102 469260
rect 511350 469248 511356 469260
rect 485096 469220 511356 469248
rect 485096 469208 485102 469220
rect 511350 469208 511356 469220
rect 511408 469208 511414 469260
rect 512638 469208 512644 469260
rect 512696 469248 512702 469260
rect 539318 469248 539324 469260
rect 512696 469220 539324 469248
rect 512696 469208 512702 469220
rect 539318 469208 539324 469220
rect 539376 469208 539382 469260
rect 540238 469208 540244 469260
rect 540296 469248 540302 469260
rect 567194 469248 567200 469260
rect 540296 469220 567200 469248
rect 540296 469208 540302 469220
rect 567194 469208 567200 469220
rect 567252 469208 567258 469260
rect 37918 468460 37924 468512
rect 37976 468500 37982 468512
rect 545758 468500 545764 468512
rect 37976 468472 545764 468500
rect 37976 468460 37982 468472
rect 545758 468460 545764 468472
rect 545816 468460 545822 468512
rect 182082 466556 182088 466608
rect 182140 466596 182146 466608
rect 233234 466596 233240 466608
rect 182140 466568 233240 466596
rect 182140 466556 182146 466568
rect 233234 466556 233240 466568
rect 233292 466556 233298 466608
rect 350442 466556 350448 466608
rect 350500 466596 350506 466608
rect 401594 466596 401600 466608
rect 350500 466568 401600 466596
rect 350500 466556 350506 466568
rect 401594 466556 401600 466568
rect 401652 466556 401658 466608
rect 462222 466556 462228 466608
rect 462280 466596 462286 466608
rect 513374 466596 513380 466608
rect 462280 466568 513380 466596
rect 462280 466556 462286 466568
rect 513374 466556 513380 466568
rect 513432 466556 513438 466608
rect 35618 466488 35624 466540
rect 35676 466528 35682 466540
rect 36814 466528 36820 466540
rect 35676 466500 36820 466528
rect 35676 466488 35682 466500
rect 36814 466488 36820 466500
rect 36872 466488 36878 466540
rect 42702 466488 42708 466540
rect 42760 466528 42766 466540
rect 93854 466528 93860 466540
rect 42760 466500 93860 466528
rect 42760 466488 42766 466500
rect 93854 466488 93860 466500
rect 93912 466488 93918 466540
rect 97902 466488 97908 466540
rect 97960 466528 97966 466540
rect 149054 466528 149060 466540
rect 97960 466500 149060 466528
rect 97960 466488 97966 466500
rect 149054 466488 149060 466500
rect 149112 466488 149118 466540
rect 154482 466488 154488 466540
rect 154540 466528 154546 466540
rect 205634 466528 205640 466540
rect 154540 466500 205640 466528
rect 154540 466488 154546 466500
rect 205634 466488 205640 466500
rect 205692 466488 205698 466540
rect 238662 466488 238668 466540
rect 238720 466528 238726 466540
rect 289814 466528 289820 466540
rect 238720 466500 289820 466528
rect 238720 466488 238726 466500
rect 289814 466488 289820 466500
rect 289872 466488 289878 466540
rect 293862 466488 293868 466540
rect 293920 466528 293926 466540
rect 345014 466528 345020 466540
rect 293920 466500 345020 466528
rect 293920 466488 293926 466500
rect 345014 466488 345020 466500
rect 345072 466488 345078 466540
rect 378042 466488 378048 466540
rect 378100 466528 378106 466540
rect 429194 466528 429200 466540
rect 378100 466500 429200 466528
rect 378100 466488 378106 466500
rect 429194 466488 429200 466500
rect 429252 466488 429258 466540
rect 434622 466488 434628 466540
rect 434680 466528 434686 466540
rect 485774 466528 485780 466540
rect 434680 466500 485780 466528
rect 434680 466488 434686 466500
rect 485774 466488 485780 466500
rect 485832 466488 485838 466540
rect 518802 466488 518808 466540
rect 518860 466528 518866 466540
rect 569954 466528 569960 466540
rect 518860 466500 569960 466528
rect 518860 466488 518866 466500
rect 569954 466488 569960 466500
rect 570012 466488 570018 466540
rect 13722 466420 13728 466472
rect 13780 466460 13786 466472
rect 66254 466460 66260 466472
rect 13780 466432 66260 466460
rect 13780 466420 13786 466432
rect 66254 466420 66260 466432
rect 66312 466420 66318 466472
rect 70302 466420 70308 466472
rect 70360 466460 70366 466472
rect 121454 466460 121460 466472
rect 70360 466432 121460 466460
rect 70360 466420 70366 466432
rect 121454 466420 121460 466432
rect 121512 466420 121518 466472
rect 126882 466420 126888 466472
rect 126940 466460 126946 466472
rect 178034 466460 178040 466472
rect 126940 466432 178040 466460
rect 126940 466420 126946 466432
rect 178034 466420 178040 466432
rect 178092 466420 178098 466472
rect 209682 466420 209688 466472
rect 209740 466460 209746 466472
rect 262214 466460 262220 466472
rect 209740 466432 262220 466460
rect 209740 466420 209746 466432
rect 262214 466420 262220 466432
rect 262272 466420 262278 466472
rect 266262 466420 266268 466472
rect 266320 466460 266326 466472
rect 317414 466460 317420 466472
rect 266320 466432 317420 466460
rect 266320 466420 266326 466432
rect 317414 466420 317420 466432
rect 317472 466420 317478 466472
rect 322842 466420 322848 466472
rect 322900 466460 322906 466472
rect 373994 466460 374000 466472
rect 322900 466432 374000 466460
rect 322900 466420 322906 466432
rect 373994 466420 374000 466432
rect 374052 466420 374058 466472
rect 405642 466420 405648 466472
rect 405700 466460 405706 466472
rect 458174 466460 458180 466472
rect 405700 466432 458180 466460
rect 405700 466420 405706 466432
rect 458174 466420 458180 466432
rect 458232 466420 458238 466472
rect 489822 466420 489828 466472
rect 489880 466460 489886 466472
rect 542354 466460 542360 466472
rect 489880 466432 542360 466460
rect 489880 466420 489886 466432
rect 542354 466420 542360 466432
rect 542412 466420 542418 466472
rect 428642 450508 428648 450560
rect 428700 450548 428706 450560
rect 435726 450548 435732 450560
rect 428700 450520 435732 450548
rect 428700 450508 428706 450520
rect 435726 450508 435732 450520
rect 435784 450508 435790 450560
rect 512730 450440 512736 450492
rect 512788 450480 512794 450492
rect 519630 450480 519636 450492
rect 512788 450452 519636 450480
rect 512788 450440 512794 450452
rect 519630 450440 519636 450452
rect 519688 450440 519694 450492
rect 483658 450304 483664 450356
rect 483716 450344 483722 450356
rect 491662 450344 491668 450356
rect 483716 450316 491668 450344
rect 483716 450304 483722 450316
rect 491662 450304 491668 450316
rect 491720 450304 491726 450356
rect 232682 449896 232688 449948
rect 232740 449936 232746 449948
rect 239766 449936 239772 449948
rect 232740 449908 239772 449936
rect 232740 449896 232746 449908
rect 239766 449896 239772 449908
rect 239824 449896 239830 449948
rect 287698 449896 287704 449948
rect 287756 449936 287762 449948
rect 295702 449936 295708 449948
rect 287756 449908 295708 449936
rect 287756 449896 287762 449908
rect 295702 449896 295708 449908
rect 295760 449896 295766 449948
rect 316770 449896 316776 449948
rect 316828 449936 316834 449948
rect 323670 449936 323676 449948
rect 316828 449908 323676 449936
rect 316828 449896 316834 449908
rect 323670 449896 323676 449908
rect 323728 449896 323734 449948
rect 63586 449624 63592 449676
rect 63644 449664 63650 449676
rect 64322 449664 64328 449676
rect 63644 449636 64328 449664
rect 63644 449624 63650 449636
rect 64322 449624 64328 449636
rect 64380 449624 64386 449676
rect 455690 449624 455696 449676
rect 455748 449664 455754 449676
rect 456150 449664 456156 449676
rect 455748 449636 456156 449664
rect 455748 449624 455754 449636
rect 456150 449624 456156 449636
rect 456208 449624 456214 449676
rect 35618 448468 35624 448520
rect 35676 448508 35682 448520
rect 36998 448508 37004 448520
rect 35676 448480 37004 448508
rect 35676 448468 35682 448480
rect 36998 448468 37004 448480
rect 37056 448468 37062 448520
rect 147674 448468 147680 448520
rect 147732 448508 147738 448520
rect 148410 448508 148416 448520
rect 147732 448480 148416 448508
rect 147732 448468 147738 448480
rect 148410 448468 148416 448480
rect 148468 448468 148474 448520
rect 343634 448468 343640 448520
rect 343692 448508 343698 448520
rect 345658 448508 345664 448520
rect 343692 448480 345664 448508
rect 343692 448468 343698 448480
rect 345658 448468 345664 448480
rect 345716 448468 345722 448520
rect 539502 448468 539508 448520
rect 539560 448508 539566 448520
rect 542998 448508 543004 448520
rect 539560 448480 543004 448508
rect 539560 448468 539566 448480
rect 542998 448468 543004 448480
rect 543056 448468 543062 448520
rect 42886 445680 42892 445732
rect 42944 445720 42950 445732
rect 72050 445720 72056 445732
rect 42944 445692 45554 445720
rect 42944 445680 42950 445692
rect 15194 445612 15200 445664
rect 15252 445652 15258 445664
rect 43990 445652 43996 445664
rect 15252 445624 43996 445652
rect 15252 445612 15258 445624
rect 43990 445612 43996 445624
rect 44048 445612 44054 445664
rect 45526 445652 45554 445692
rect 64846 445692 72056 445720
rect 64846 445652 64874 445692
rect 72050 445680 72056 445692
rect 72108 445680 72114 445732
rect 99466 445680 99472 445732
rect 99524 445720 99530 445732
rect 99524 445692 103514 445720
rect 99524 445680 99530 445692
rect 45526 445624 64874 445652
rect 71866 445612 71872 445664
rect 71924 445652 71930 445664
rect 100018 445652 100024 445664
rect 71924 445624 100024 445652
rect 71924 445612 71930 445624
rect 100018 445612 100024 445624
rect 100076 445612 100082 445664
rect 103486 445652 103514 445692
rect 127066 445680 127072 445732
rect 127124 445720 127130 445732
rect 127124 445692 132494 445720
rect 127124 445680 127130 445692
rect 127986 445652 127992 445664
rect 103486 445624 127992 445652
rect 127986 445612 127992 445624
rect 128044 445612 128050 445664
rect 132466 445652 132494 445692
rect 183646 445680 183652 445732
rect 183704 445720 183710 445732
rect 183704 445692 190454 445720
rect 183704 445680 183710 445692
rect 156046 445652 156052 445664
rect 132466 445624 156052 445652
rect 156046 445612 156052 445624
rect 156104 445612 156110 445664
rect 165982 445612 165988 445664
rect 166040 445652 166046 445664
rect 177298 445652 177304 445664
rect 166040 445624 177304 445652
rect 166040 445612 166046 445624
rect 177298 445612 177304 445624
rect 177356 445612 177362 445664
rect 178678 445612 178684 445664
rect 178736 445652 178742 445664
rect 184014 445652 184020 445664
rect 178736 445624 184020 445652
rect 178736 445612 178742 445624
rect 184014 445612 184020 445624
rect 184072 445612 184078 445664
rect 190426 445652 190454 445692
rect 374638 445680 374644 445732
rect 374696 445720 374702 445732
rect 379698 445720 379704 445732
rect 374696 445692 379704 445720
rect 374696 445680 374702 445692
rect 379698 445680 379704 445692
rect 379756 445680 379762 445732
rect 211706 445652 211712 445664
rect 190426 445624 211712 445652
rect 211706 445612 211712 445624
rect 211764 445612 211770 445664
rect 222010 445612 222016 445664
rect 222068 445652 222074 445664
rect 232590 445652 232596 445664
rect 222068 445624 232596 445652
rect 222068 445612 222074 445624
rect 232590 445612 232596 445624
rect 232648 445612 232654 445664
rect 249702 445612 249708 445664
rect 249760 445652 249766 445664
rect 260190 445652 260196 445664
rect 249760 445624 260196 445652
rect 249760 445612 249766 445624
rect 260190 445612 260196 445624
rect 260248 445612 260254 445664
rect 261478 445612 261484 445664
rect 261536 445652 261542 445664
rect 567194 445652 567200 445664
rect 261536 445624 567200 445652
rect 261536 445612 261542 445624
rect 567194 445612 567200 445624
rect 567252 445612 567258 445664
rect 25682 445544 25688 445596
rect 25740 445584 25746 445596
rect 36906 445584 36912 445596
rect 25740 445556 36912 445584
rect 25740 445544 25746 445556
rect 36906 445544 36912 445556
rect 36964 445544 36970 445596
rect 53650 445544 53656 445596
rect 53708 445584 53714 445596
rect 69658 445584 69664 445596
rect 53708 445556 69664 445584
rect 53708 445544 53714 445556
rect 69658 445544 69664 445556
rect 69716 445544 69722 445596
rect 81986 445544 81992 445596
rect 82044 445584 82050 445596
rect 94498 445584 94504 445596
rect 82044 445556 94504 445584
rect 82044 445544 82050 445556
rect 94498 445544 94504 445556
rect 94556 445544 94562 445596
rect 109678 445544 109684 445596
rect 109736 445584 109742 445596
rect 120718 445584 120724 445596
rect 109736 445556 120724 445584
rect 109736 445544 109742 445556
rect 120718 445544 120724 445556
rect 120776 445544 120782 445596
rect 137646 445544 137652 445596
rect 137704 445584 137710 445596
rect 148318 445584 148324 445596
rect 137704 445556 148324 445584
rect 137704 445544 137710 445556
rect 148318 445544 148324 445556
rect 148376 445544 148382 445596
rect 193674 445544 193680 445596
rect 193732 445584 193738 445596
rect 204898 445584 204904 445596
rect 193732 445556 204904 445584
rect 193732 445544 193738 445556
rect 204898 445544 204904 445556
rect 204956 445544 204962 445596
rect 238846 445544 238852 445596
rect 238904 445584 238910 445596
rect 268010 445584 268016 445596
rect 238904 445556 268016 445584
rect 238904 445544 238910 445556
rect 268010 445544 268016 445556
rect 268068 445544 268074 445596
rect 277670 445544 277676 445596
rect 277728 445584 277734 445596
rect 289078 445584 289084 445596
rect 277728 445556 289084 445584
rect 277728 445544 277734 445556
rect 289078 445544 289084 445556
rect 289136 445544 289142 445596
rect 306006 445544 306012 445596
rect 306064 445584 306070 445596
rect 316678 445584 316684 445596
rect 306064 445556 316684 445584
rect 306064 445544 306070 445556
rect 316678 445544 316684 445556
rect 316736 445544 316742 445596
rect 323026 445544 323032 445596
rect 323084 445584 323090 445596
rect 352006 445584 352012 445596
rect 323084 445556 352012 445584
rect 323084 445544 323090 445556
rect 352006 445544 352012 445556
rect 352064 445544 352070 445596
rect 361666 445544 361672 445596
rect 361724 445584 361730 445596
rect 373258 445584 373264 445596
rect 361724 445556 373264 445584
rect 361724 445544 361730 445556
rect 373258 445544 373264 445556
rect 373316 445544 373322 445596
rect 379606 445544 379612 445596
rect 379664 445584 379670 445596
rect 408034 445584 408040 445596
rect 379664 445556 408040 445584
rect 379664 445544 379670 445556
rect 408034 445544 408040 445556
rect 408092 445544 408098 445596
rect 417694 445544 417700 445596
rect 417752 445584 417758 445596
rect 428550 445584 428556 445596
rect 417752 445556 428556 445584
rect 417752 445544 417758 445556
rect 428550 445544 428556 445556
rect 428608 445544 428614 445596
rect 434806 445544 434812 445596
rect 434864 445584 434870 445596
rect 463694 445584 463700 445596
rect 434864 445556 463700 445584
rect 434864 445544 434870 445556
rect 463694 445544 463700 445556
rect 463752 445544 463758 445596
rect 473998 445544 474004 445596
rect 474056 445584 474062 445596
rect 485038 445584 485044 445596
rect 474056 445556 485044 445584
rect 474056 445544 474062 445556
rect 485038 445544 485044 445556
rect 485096 445544 485102 445596
rect 501690 445544 501696 445596
rect 501748 445584 501754 445596
rect 512638 445584 512644 445596
rect 501748 445556 512644 445584
rect 501748 445544 501754 445556
rect 512638 445544 512644 445556
rect 512696 445544 512702 445596
rect 518986 445544 518992 445596
rect 519044 445584 519050 445596
rect 547874 445584 547880 445596
rect 519044 445556 547880 445584
rect 519044 445544 519050 445556
rect 547874 445544 547880 445556
rect 547932 445544 547938 445596
rect 333698 445476 333704 445528
rect 333756 445516 333762 445528
rect 344278 445516 344284 445528
rect 333756 445488 344284 445516
rect 333756 445476 333762 445488
rect 344278 445476 344284 445488
rect 344336 445476 344342 445528
rect 390002 445476 390008 445528
rect 390060 445516 390066 445528
rect 400858 445516 400864 445528
rect 390060 445488 400864 445516
rect 390060 445476 390066 445488
rect 400858 445476 400864 445488
rect 400916 445476 400922 445528
rect 445662 445476 445668 445528
rect 445720 445516 445726 445528
rect 456058 445516 456064 445528
rect 445720 445488 456064 445516
rect 445720 445476 445726 445488
rect 456058 445476 456064 445488
rect 456116 445476 456122 445528
rect 529658 445476 529664 445528
rect 529716 445516 529722 445528
rect 540238 445516 540244 445528
rect 529716 445488 540244 445516
rect 529716 445476 529722 445488
rect 540238 445476 540244 445488
rect 540296 445476 540302 445528
rect 36722 445408 36728 445460
rect 36780 445448 36786 445460
rect 557534 445448 557540 445460
rect 36780 445420 557540 445448
rect 36780 445408 36786 445420
rect 557534 445408 557540 445420
rect 557592 445408 557598 445460
rect 16022 443640 16028 443692
rect 16080 443680 16086 443692
rect 547874 443680 547880 443692
rect 16080 443652 547880 443680
rect 16080 443640 16086 443652
rect 547874 443640 547880 443652
rect 547932 443640 547938 443692
rect 25682 443164 25688 443216
rect 25740 443204 25746 443216
rect 69658 443204 69664 443216
rect 25740 443176 69664 443204
rect 25740 443164 25746 443176
rect 69658 443164 69664 443176
rect 69716 443164 69722 443216
rect 212258 443164 212264 443216
rect 212316 443204 212322 443216
rect 232682 443204 232688 443216
rect 212316 443176 232688 443204
rect 212316 443164 212322 443176
rect 232682 443164 232688 443176
rect 232740 443164 232746 443216
rect 296346 443164 296352 443216
rect 296404 443204 296410 443216
rect 316770 443204 316776 443216
rect 296404 443176 316776 443204
rect 296404 443164 296410 443176
rect 316770 443164 316776 443176
rect 316828 443164 316834 443216
rect 408034 443164 408040 443216
rect 408092 443204 408098 443216
rect 428642 443204 428648 443216
rect 408092 443176 428648 443204
rect 408092 443164 408098 443176
rect 428642 443164 428648 443176
rect 428700 443164 428706 443216
rect 492030 443164 492036 443216
rect 492088 443204 492094 443216
rect 512730 443204 512736 443216
rect 492088 443176 512736 443204
rect 492088 443164 492094 443176
rect 512730 443164 512736 443176
rect 512788 443164 512794 443216
rect 36906 443096 36912 443148
rect 36964 443136 36970 443148
rect 53374 443136 53380 443148
rect 36964 443108 53380 443136
rect 36964 443096 36970 443108
rect 53374 443096 53380 443108
rect 53432 443096 53438 443148
rect 64322 443096 64328 443148
rect 64380 443136 64386 443148
rect 81434 443136 81440 443148
rect 64380 443108 81440 443136
rect 64380 443096 64386 443108
rect 81434 443096 81440 443108
rect 81492 443096 81498 443148
rect 148318 443096 148324 443148
rect 148376 443136 148382 443148
rect 165614 443136 165620 443148
rect 148376 443108 165620 443136
rect 148376 443096 148382 443108
rect 165614 443096 165620 443108
rect 165672 443096 165678 443148
rect 175458 443096 175464 443148
rect 175516 443136 175522 443148
rect 193674 443136 193680 443148
rect 175516 443108 193680 443136
rect 175516 443096 175522 443108
rect 193674 443096 193680 443108
rect 193732 443096 193738 443148
rect 203518 443096 203524 443148
rect 203576 443136 203582 443148
rect 221366 443136 221372 443148
rect 203576 443108 221372 443136
rect 203576 443096 203582 443108
rect 221366 443096 221372 443108
rect 221424 443096 221430 443148
rect 260190 443096 260196 443148
rect 260248 443136 260254 443148
rect 277670 443136 277676 443148
rect 260248 443108 277676 443136
rect 260248 443096 260254 443108
rect 277670 443096 277676 443108
rect 277728 443096 277734 443148
rect 287514 443096 287520 443148
rect 287572 443136 287578 443148
rect 305362 443136 305368 443148
rect 287572 443108 305368 443136
rect 287572 443096 287578 443108
rect 305362 443096 305368 443108
rect 305420 443096 305426 443148
rect 345658 443096 345664 443148
rect 345716 443136 345722 443148
rect 361666 443136 361672 443148
rect 345716 443108 361672 443136
rect 345716 443096 345722 443108
rect 361666 443096 361672 443108
rect 361724 443096 361730 443148
rect 371510 443096 371516 443148
rect 371568 443136 371574 443148
rect 389358 443136 389364 443148
rect 371568 443108 389364 443136
rect 371568 443096 371574 443108
rect 389358 443096 389364 443108
rect 389416 443096 389422 443148
rect 399478 443096 399484 443148
rect 399536 443136 399542 443148
rect 417694 443136 417700 443148
rect 399536 443108 417700 443136
rect 399536 443096 399542 443108
rect 417694 443096 417700 443108
rect 417752 443096 417758 443148
rect 456058 443096 456064 443148
rect 456116 443136 456122 443148
rect 473538 443136 473544 443148
rect 456116 443108 473544 443136
rect 456116 443096 456122 443108
rect 473538 443096 473544 443108
rect 473596 443096 473602 443148
rect 483474 443096 483480 443148
rect 483532 443136 483538 443148
rect 501690 443136 501696 443148
rect 483532 443108 501696 443136
rect 483532 443096 483538 443108
rect 501690 443096 501696 443108
rect 501748 443096 501754 443148
rect 36998 443028 37004 443080
rect 37056 443068 37062 443080
rect 62942 443068 62948 443080
rect 37056 443040 62948 443068
rect 37056 443028 37062 443040
rect 62942 443028 62948 443040
rect 63000 443028 63006 443080
rect 66898 443028 66904 443080
rect 66956 443068 66962 443080
rect 91094 443068 91100 443080
rect 66956 443040 91100 443068
rect 66956 443028 66962 443040
rect 91094 443028 91100 443040
rect 91152 443028 91158 443080
rect 91462 443028 91468 443080
rect 91520 443068 91526 443080
rect 109678 443068 109684 443080
rect 91520 443040 109684 443068
rect 91520 443028 91526 443040
rect 109678 443028 109684 443040
rect 109736 443028 109742 443080
rect 119430 443028 119436 443080
rect 119488 443068 119494 443080
rect 137278 443068 137284 443080
rect 119488 443040 137284 443068
rect 119488 443028 119494 443040
rect 137278 443028 137284 443040
rect 137336 443028 137342 443080
rect 156322 443028 156328 443080
rect 156380 443068 156386 443080
rect 178678 443068 178684 443080
rect 156380 443040 178684 443068
rect 156380 443028 156386 443040
rect 178678 443028 178684 443040
rect 178736 443028 178742 443080
rect 232498 443028 232504 443080
rect 232556 443068 232562 443080
rect 249334 443068 249340 443080
rect 232556 443040 249340 443068
rect 232556 443028 232562 443040
rect 249334 443028 249340 443040
rect 249392 443028 249398 443080
rect 268010 443028 268016 443080
rect 268068 443068 268074 443080
rect 287698 443068 287704 443080
rect 268068 443040 287704 443068
rect 268068 443028 268074 443040
rect 287698 443028 287704 443040
rect 287756 443028 287762 443080
rect 315482 443028 315488 443080
rect 315540 443068 315546 443080
rect 333422 443068 333428 443080
rect 315540 443040 333428 443068
rect 315540 443028 315546 443040
rect 333422 443028 333428 443040
rect 333480 443028 333486 443080
rect 352006 443028 352012 443080
rect 352064 443068 352070 443080
rect 374638 443068 374644 443080
rect 352064 443040 374644 443068
rect 352064 443028 352070 443040
rect 374638 443028 374644 443040
rect 374696 443028 374702 443080
rect 428550 443028 428556 443080
rect 428608 443068 428614 443080
rect 445662 443068 445668 443080
rect 428608 443040 445668 443068
rect 428608 443028 428614 443040
rect 445662 443028 445668 443040
rect 445720 443028 445726 443080
rect 464338 443028 464344 443080
rect 464396 443068 464402 443080
rect 483658 443068 483664 443080
rect 464396 443040 483664 443068
rect 464396 443028 464402 443040
rect 483658 443028 483664 443040
rect 483716 443028 483722 443080
rect 511442 443028 511448 443080
rect 511500 443068 511506 443080
rect 529658 443068 529664 443080
rect 511500 443040 529664 443068
rect 511500 443028 511506 443040
rect 529658 443028 529664 443040
rect 529716 443028 529722 443080
rect 542998 443028 543004 443080
rect 543056 443068 543062 443080
rect 557534 443068 557540 443080
rect 543056 443040 557540 443068
rect 543056 443028 543062 443040
rect 557534 443028 557540 443040
rect 557592 443028 557598 443080
rect 94498 442960 94504 443012
rect 94556 443000 94562 443012
rect 119338 443000 119344 443012
rect 94556 442972 119344 443000
rect 94556 442960 94562 442972
rect 119338 442960 119344 442972
rect 119396 442960 119402 443012
rect 120718 442960 120724 443012
rect 120776 443000 120782 443012
rect 147030 443000 147036 443012
rect 120776 442972 147036 443000
rect 120776 442960 120782 442972
rect 147030 442960 147036 442972
rect 147088 442960 147094 443012
rect 148410 442960 148416 443012
rect 148468 443000 148474 443012
rect 175274 443000 175280 443012
rect 148468 442972 175280 443000
rect 148468 442960 148474 442972
rect 175274 442960 175280 442972
rect 175332 442960 175338 443012
rect 177298 442960 177304 443012
rect 177356 443000 177362 443012
rect 203334 443000 203340 443012
rect 177356 442972 203340 443000
rect 177356 442960 177362 442972
rect 203334 442960 203340 442972
rect 203392 442960 203398 443012
rect 204898 442960 204904 443012
rect 204956 443000 204962 443012
rect 231026 443000 231032 443012
rect 204956 442972 231032 443000
rect 204956 442960 204962 442972
rect 231026 442960 231032 442972
rect 231084 442960 231090 443012
rect 232590 442960 232596 443012
rect 232648 443000 232654 443012
rect 259086 443000 259092 443012
rect 232648 442972 259092 443000
rect 232648 442960 232654 442972
rect 259086 442960 259092 442972
rect 259144 442960 259150 443012
rect 260098 442960 260104 443012
rect 260156 443000 260162 443012
rect 287330 443000 287336 443012
rect 260156 442972 287336 443000
rect 260156 442960 260162 442972
rect 287330 442960 287336 442972
rect 287388 442960 287394 443012
rect 289078 442960 289084 443012
rect 289136 443000 289142 443012
rect 315022 443000 315028 443012
rect 289136 442972 315028 443000
rect 289136 442960 289142 442972
rect 315022 442960 315028 442972
rect 315080 442960 315086 443012
rect 316678 442960 316684 443012
rect 316736 443000 316742 443012
rect 342990 443000 342996 443012
rect 316736 442972 342996 443000
rect 316736 442960 316742 442972
rect 342990 442960 342996 442972
rect 343048 442960 343054 443012
rect 344278 442960 344284 443012
rect 344336 443000 344342 443012
rect 371326 443000 371332 443012
rect 344336 442972 371332 443000
rect 344336 442960 344342 442972
rect 371326 442960 371332 442972
rect 371384 442960 371390 443012
rect 373258 442960 373264 443012
rect 373316 443000 373322 443012
rect 399018 443000 399024 443012
rect 373316 442972 399024 443000
rect 373316 442960 373322 442972
rect 399018 442960 399024 442972
rect 399076 442960 399082 443012
rect 400858 442960 400864 443012
rect 400916 443000 400922 443012
rect 427354 443000 427360 443012
rect 400916 442972 427360 443000
rect 400916 442960 400922 442972
rect 427354 442960 427360 442972
rect 427412 442960 427418 443012
rect 428458 442960 428464 443012
rect 428516 443000 428522 443012
rect 455322 443000 455328 443012
rect 428516 442972 455328 443000
rect 428516 442960 428522 442972
rect 455322 442960 455328 442972
rect 455380 442960 455386 443012
rect 456150 442960 456156 443012
rect 456208 443000 456214 443012
rect 483198 443000 483204 443012
rect 456208 442972 483204 443000
rect 456208 442960 456214 442972
rect 483198 442960 483204 442972
rect 483256 442960 483262 443012
rect 485038 442960 485044 443012
rect 485096 443000 485102 443012
rect 511350 443000 511356 443012
rect 485096 442972 511356 443000
rect 485096 442960 485102 442972
rect 511350 442960 511356 442972
rect 511408 442960 511414 443012
rect 512638 442960 512644 443012
rect 512696 443000 512702 443012
rect 539318 443000 539324 443012
rect 512696 442972 539324 443000
rect 512696 442960 512702 442972
rect 539318 442960 539324 442972
rect 539376 442960 539382 443012
rect 540238 442960 540244 443012
rect 540296 443000 540302 443012
rect 567194 443000 567200 443012
rect 540296 442972 567200 443000
rect 540296 442960 540302 442972
rect 567194 442960 567200 442972
rect 567252 442960 567258 443012
rect 37918 440852 37924 440904
rect 37976 440892 37982 440904
rect 545758 440892 545764 440904
rect 37976 440864 545764 440892
rect 37976 440852 37982 440864
rect 545758 440852 545764 440864
rect 545816 440852 545822 440904
rect 182082 440308 182088 440360
rect 182140 440348 182146 440360
rect 233234 440348 233240 440360
rect 182140 440320 233240 440348
rect 182140 440308 182146 440320
rect 233234 440308 233240 440320
rect 233292 440308 233298 440360
rect 350442 440308 350448 440360
rect 350500 440348 350506 440360
rect 401594 440348 401600 440360
rect 350500 440320 401600 440348
rect 350500 440308 350506 440320
rect 401594 440308 401600 440320
rect 401652 440308 401658 440360
rect 35618 440240 35624 440292
rect 35676 440280 35682 440292
rect 36722 440280 36728 440292
rect 35676 440252 36728 440280
rect 35676 440240 35682 440252
rect 36722 440240 36728 440252
rect 36780 440240 36786 440292
rect 42702 440240 42708 440292
rect 42760 440280 42766 440292
rect 93854 440280 93860 440292
rect 42760 440252 93860 440280
rect 42760 440240 42766 440252
rect 93854 440240 93860 440252
rect 93912 440240 93918 440292
rect 97902 440240 97908 440292
rect 97960 440280 97966 440292
rect 149054 440280 149060 440292
rect 97960 440252 149060 440280
rect 97960 440240 97966 440252
rect 149054 440240 149060 440252
rect 149112 440240 149118 440292
rect 154482 440240 154488 440292
rect 154540 440280 154546 440292
rect 205634 440280 205640 440292
rect 154540 440252 205640 440280
rect 154540 440240 154546 440252
rect 205634 440240 205640 440252
rect 205692 440240 205698 440292
rect 238662 440240 238668 440292
rect 238720 440280 238726 440292
rect 289814 440280 289820 440292
rect 238720 440252 289820 440280
rect 238720 440240 238726 440252
rect 289814 440240 289820 440252
rect 289872 440240 289878 440292
rect 293862 440240 293868 440292
rect 293920 440280 293926 440292
rect 345014 440280 345020 440292
rect 293920 440252 345020 440280
rect 293920 440240 293926 440252
rect 345014 440240 345020 440252
rect 345072 440240 345078 440292
rect 378042 440240 378048 440292
rect 378100 440280 378106 440292
rect 429194 440280 429200 440292
rect 378100 440252 429200 440280
rect 378100 440240 378106 440252
rect 429194 440240 429200 440252
rect 429252 440240 429258 440292
rect 434622 440240 434628 440292
rect 434680 440280 434686 440292
rect 485774 440280 485780 440292
rect 434680 440252 485780 440280
rect 434680 440240 434686 440252
rect 485774 440240 485780 440252
rect 485832 440240 485838 440292
rect 489822 440240 489828 440292
rect 489880 440280 489886 440292
rect 542354 440280 542360 440292
rect 489880 440252 542360 440280
rect 489880 440240 489886 440252
rect 542354 440240 542360 440252
rect 542412 440240 542418 440292
rect 63586 427116 63592 427168
rect 63644 427156 63650 427168
rect 64322 427156 64328 427168
rect 63644 427128 64328 427156
rect 63644 427116 63650 427128
rect 64322 427116 64328 427128
rect 64380 427116 64386 427168
rect 259730 427116 259736 427168
rect 259788 427156 259794 427168
rect 260190 427156 260196 427168
rect 259788 427128 260196 427156
rect 259788 427116 259794 427128
rect 260190 427116 260196 427128
rect 260248 427116 260254 427168
rect 287698 423580 287704 423632
rect 287756 423620 287762 423632
rect 295702 423620 295708 423632
rect 287756 423592 295708 423620
rect 287756 423580 287762 423592
rect 295702 423580 295708 423592
rect 295760 423580 295766 423632
rect 316770 423580 316776 423632
rect 316828 423620 316834 423632
rect 323670 423620 323676 423632
rect 316828 423592 323676 423620
rect 316828 423580 316834 423592
rect 323670 423580 323676 423592
rect 323728 423580 323734 423632
rect 483658 423036 483664 423088
rect 483716 423076 483722 423088
rect 491662 423076 491668 423088
rect 483716 423048 491668 423076
rect 483716 423036 483722 423048
rect 491662 423036 491668 423048
rect 491720 423036 491726 423088
rect 232682 422968 232688 423020
rect 232740 423008 232746 423020
rect 239766 423008 239772 423020
rect 232740 422980 239772 423008
rect 232740 422968 232746 422980
rect 239766 422968 239772 422980
rect 239824 422968 239830 423020
rect 512730 422968 512736 423020
rect 512788 423008 512794 423020
rect 519630 423008 519636 423020
rect 512788 422980 519636 423008
rect 512788 422968 512794 422980
rect 519630 422968 519636 422980
rect 519688 422968 519694 423020
rect 428642 422900 428648 422952
rect 428700 422940 428706 422952
rect 435726 422940 435732 422952
rect 428700 422912 435732 422940
rect 428700 422900 428706 422912
rect 435726 422900 435732 422912
rect 435784 422900 435790 422952
rect 13722 422220 13728 422272
rect 13780 422260 13786 422272
rect 66254 422260 66260 422272
rect 13780 422232 66260 422260
rect 13780 422220 13786 422232
rect 66254 422220 66260 422232
rect 66312 422220 66318 422272
rect 70302 422220 70308 422272
rect 70360 422260 70366 422272
rect 121454 422260 121460 422272
rect 70360 422232 121460 422260
rect 70360 422220 70366 422232
rect 121454 422220 121460 422232
rect 121512 422220 121518 422272
rect 126882 422220 126888 422272
rect 126940 422260 126946 422272
rect 178034 422260 178040 422272
rect 126940 422232 178040 422260
rect 126940 422220 126946 422232
rect 178034 422220 178040 422232
rect 178092 422220 178098 422272
rect 209682 422220 209688 422272
rect 209740 422260 209746 422272
rect 262214 422260 262220 422272
rect 209740 422232 262220 422260
rect 209740 422220 209746 422232
rect 262214 422220 262220 422232
rect 262272 422220 262278 422272
rect 266262 422220 266268 422272
rect 266320 422260 266326 422272
rect 317414 422260 317420 422272
rect 266320 422232 317420 422260
rect 266320 422220 266326 422232
rect 317414 422220 317420 422232
rect 317472 422220 317478 422272
rect 322842 422220 322848 422272
rect 322900 422260 322906 422272
rect 373994 422260 374000 422272
rect 322900 422232 374000 422260
rect 322900 422220 322906 422232
rect 373994 422220 374000 422232
rect 374052 422220 374058 422272
rect 405642 422220 405648 422272
rect 405700 422260 405706 422272
rect 458174 422260 458180 422272
rect 405700 422232 458180 422260
rect 405700 422220 405706 422232
rect 458174 422220 458180 422232
rect 458232 422220 458238 422272
rect 462222 422220 462228 422272
rect 462280 422260 462286 422272
rect 513374 422260 513380 422272
rect 462280 422232 513380 422260
rect 462280 422220 462286 422232
rect 513374 422220 513380 422232
rect 513432 422220 513438 422272
rect 518802 422220 518808 422272
rect 518860 422260 518866 422272
rect 569954 422260 569960 422272
rect 518860 422232 569960 422260
rect 518860 422220 518866 422232
rect 569954 422220 569960 422232
rect 570012 422220 570018 422272
rect 35618 422152 35624 422204
rect 35676 422192 35682 422204
rect 36906 422192 36912 422204
rect 35676 422164 36912 422192
rect 35676 422152 35682 422164
rect 36906 422152 36912 422164
rect 36964 422152 36970 422204
rect 343542 422152 343548 422204
rect 343600 422192 343606 422204
rect 345658 422192 345664 422204
rect 343600 422164 345664 422192
rect 343600 422152 343606 422164
rect 345658 422152 345664 422164
rect 345716 422152 345722 422204
rect 427722 421676 427728 421728
rect 427780 421716 427786 421728
rect 428550 421716 428556 421728
rect 427780 421688 428556 421716
rect 427780 421676 427786 421688
rect 428550 421676 428556 421688
rect 428608 421676 428614 421728
rect 539502 421676 539508 421728
rect 539560 421716 539566 421728
rect 542998 421716 543004 421728
rect 539560 421688 543004 421716
rect 539560 421676 539566 421688
rect 542998 421676 543004 421688
rect 543056 421676 543062 421728
rect 178678 419432 178684 419484
rect 178736 419472 178742 419484
rect 184014 419472 184020 419484
rect 178736 419444 184020 419472
rect 178736 419432 178742 419444
rect 184014 419432 184020 419444
rect 184072 419432 184078 419484
rect 374638 419432 374644 419484
rect 374696 419472 374702 419484
rect 379698 419472 379704 419484
rect 374696 419444 379704 419472
rect 374696 419432 374702 419444
rect 379698 419432 379704 419444
rect 379756 419432 379762 419484
rect 15194 419364 15200 419416
rect 15252 419404 15258 419416
rect 43990 419404 43996 419416
rect 15252 419376 43996 419404
rect 15252 419364 15258 419376
rect 43990 419364 43996 419376
rect 44048 419364 44054 419416
rect 71038 419364 71044 419416
rect 71096 419404 71102 419416
rect 567194 419404 567200 419416
rect 71096 419376 567200 419404
rect 71096 419364 71102 419376
rect 567194 419364 567200 419376
rect 567252 419364 567258 419416
rect 25682 419296 25688 419348
rect 25740 419336 25746 419348
rect 36998 419336 37004 419348
rect 25740 419308 37004 419336
rect 25740 419296 25746 419308
rect 36998 419296 37004 419308
rect 37056 419296 37062 419348
rect 53650 419296 53656 419348
rect 53708 419336 53714 419348
rect 66898 419336 66904 419348
rect 53708 419308 66904 419336
rect 53708 419296 53714 419308
rect 66898 419296 66904 419308
rect 66956 419296 66962 419348
rect 71866 419296 71872 419348
rect 71924 419336 71930 419348
rect 100018 419336 100024 419348
rect 71924 419308 100024 419336
rect 71924 419296 71930 419308
rect 100018 419296 100024 419308
rect 100076 419296 100082 419348
rect 127986 419336 127992 419348
rect 103486 419308 127992 419336
rect 42886 419228 42892 419280
rect 42944 419268 42950 419280
rect 72050 419268 72056 419280
rect 42944 419240 72056 419268
rect 42944 419228 42950 419240
rect 72050 419228 72056 419240
rect 72108 419228 72114 419280
rect 81986 419228 81992 419280
rect 82044 419268 82050 419280
rect 94498 419268 94504 419280
rect 82044 419240 94504 419268
rect 82044 419228 82050 419240
rect 94498 419228 94504 419240
rect 94556 419228 94562 419280
rect 99466 419228 99472 419280
rect 99524 419268 99530 419280
rect 103486 419268 103514 419308
rect 127986 419296 127992 419308
rect 128044 419296 128050 419348
rect 156046 419336 156052 419348
rect 132466 419308 156052 419336
rect 99524 419240 103514 419268
rect 99524 419228 99530 419240
rect 109678 419228 109684 419280
rect 109736 419268 109742 419280
rect 120718 419268 120724 419280
rect 109736 419240 120724 419268
rect 109736 419228 109742 419240
rect 120718 419228 120724 419240
rect 120776 419228 120782 419280
rect 127066 419228 127072 419280
rect 127124 419268 127130 419280
rect 132466 419268 132494 419308
rect 156046 419296 156052 419308
rect 156104 419296 156110 419348
rect 165982 419296 165988 419348
rect 166040 419336 166046 419348
rect 177298 419336 177304 419348
rect 166040 419308 177304 419336
rect 166040 419296 166046 419308
rect 177298 419296 177304 419308
rect 177356 419296 177362 419348
rect 183646 419296 183652 419348
rect 183704 419336 183710 419348
rect 211706 419336 211712 419348
rect 183704 419308 211712 419336
rect 183704 419296 183710 419308
rect 211706 419296 211712 419308
rect 211764 419296 211770 419348
rect 222010 419296 222016 419348
rect 222068 419336 222074 419348
rect 232590 419336 232596 419348
rect 222068 419308 232596 419336
rect 222068 419296 222074 419308
rect 232590 419296 232596 419308
rect 232648 419296 232654 419348
rect 238846 419296 238852 419348
rect 238904 419336 238910 419348
rect 268010 419336 268016 419348
rect 238904 419308 268016 419336
rect 238904 419296 238910 419308
rect 268010 419296 268016 419308
rect 268068 419296 268074 419348
rect 277670 419296 277676 419348
rect 277728 419336 277734 419348
rect 289078 419336 289084 419348
rect 277728 419308 289084 419336
rect 277728 419296 277734 419308
rect 289078 419296 289084 419308
rect 289136 419296 289142 419348
rect 306006 419296 306012 419348
rect 306064 419336 306070 419348
rect 316678 419336 316684 419348
rect 306064 419308 316684 419336
rect 306064 419296 306070 419308
rect 316678 419296 316684 419308
rect 316736 419296 316742 419348
rect 323026 419296 323032 419348
rect 323084 419336 323090 419348
rect 352006 419336 352012 419348
rect 323084 419308 352012 419336
rect 323084 419296 323090 419308
rect 352006 419296 352012 419308
rect 352064 419296 352070 419348
rect 361666 419296 361672 419348
rect 361724 419336 361730 419348
rect 373258 419336 373264 419348
rect 361724 419308 373264 419336
rect 361724 419296 361730 419308
rect 373258 419296 373264 419308
rect 373316 419296 373322 419348
rect 379606 419296 379612 419348
rect 379664 419336 379670 419348
rect 408034 419336 408040 419348
rect 379664 419308 408040 419336
rect 379664 419296 379670 419308
rect 408034 419296 408040 419308
rect 408092 419296 408098 419348
rect 417694 419296 417700 419348
rect 417752 419336 417758 419348
rect 428458 419336 428464 419348
rect 417752 419308 428464 419336
rect 417752 419296 417758 419308
rect 428458 419296 428464 419308
rect 428516 419296 428522 419348
rect 434806 419296 434812 419348
rect 434864 419336 434870 419348
rect 463694 419336 463700 419348
rect 434864 419308 463700 419336
rect 434864 419296 434870 419308
rect 463694 419296 463700 419308
rect 463752 419296 463758 419348
rect 473998 419296 474004 419348
rect 474056 419336 474062 419348
rect 485038 419336 485044 419348
rect 474056 419308 485044 419336
rect 474056 419296 474062 419308
rect 485038 419296 485044 419308
rect 485096 419296 485102 419348
rect 501690 419296 501696 419348
rect 501748 419336 501754 419348
rect 512638 419336 512644 419348
rect 501748 419308 512644 419336
rect 501748 419296 501754 419308
rect 512638 419296 512644 419308
rect 512696 419296 512702 419348
rect 518986 419296 518992 419348
rect 519044 419336 519050 419348
rect 547874 419336 547880 419348
rect 519044 419308 547880 419336
rect 519044 419296 519050 419308
rect 547874 419296 547880 419308
rect 547932 419296 547938 419348
rect 127124 419240 132494 419268
rect 127124 419228 127130 419240
rect 137646 419228 137652 419280
rect 137704 419268 137710 419280
rect 148410 419268 148416 419280
rect 137704 419240 148416 419268
rect 137704 419228 137710 419240
rect 148410 419228 148416 419240
rect 148468 419228 148474 419280
rect 193674 419228 193680 419280
rect 193732 419268 193738 419280
rect 204898 419268 204904 419280
rect 193732 419240 204904 419268
rect 193732 419228 193738 419240
rect 204898 419228 204904 419240
rect 204956 419228 204962 419280
rect 249702 419228 249708 419280
rect 249760 419268 249766 419280
rect 260098 419268 260104 419280
rect 249760 419240 260104 419268
rect 249760 419228 249766 419240
rect 260098 419228 260104 419240
rect 260156 419228 260162 419280
rect 333698 419228 333704 419280
rect 333756 419268 333762 419280
rect 344278 419268 344284 419280
rect 333756 419240 344284 419268
rect 333756 419228 333762 419240
rect 344278 419228 344284 419240
rect 344336 419228 344342 419280
rect 390002 419228 390008 419280
rect 390060 419268 390066 419280
rect 400858 419268 400864 419280
rect 390060 419240 400864 419268
rect 390060 419228 390066 419240
rect 400858 419228 400864 419240
rect 400916 419228 400922 419280
rect 445662 419228 445668 419280
rect 445720 419268 445726 419280
rect 456150 419268 456156 419280
rect 445720 419240 456156 419268
rect 445720 419228 445726 419240
rect 456150 419228 456156 419240
rect 456208 419228 456214 419280
rect 529658 419228 529664 419280
rect 529716 419268 529722 419280
rect 540238 419268 540244 419280
rect 529716 419240 540244 419268
rect 529716 419228 529722 419240
rect 540238 419228 540244 419240
rect 540296 419228 540302 419280
rect 36814 419160 36820 419212
rect 36872 419200 36878 419212
rect 557534 419200 557540 419212
rect 36872 419172 557540 419200
rect 36872 419160 36878 419172
rect 557534 419160 557540 419172
rect 557592 419160 557598 419212
rect 16022 416032 16028 416084
rect 16080 416072 16086 416084
rect 547874 416072 547880 416084
rect 16080 416044 547880 416072
rect 16080 416032 16086 416044
rect 547874 416032 547880 416044
rect 547932 416032 547938 416084
rect 25682 415692 25688 415744
rect 25740 415732 25746 415744
rect 261478 415732 261484 415744
rect 25740 415704 261484 415732
rect 25740 415692 25746 415704
rect 261478 415692 261484 415704
rect 261536 415692 261542 415744
rect 119430 415624 119436 415676
rect 119488 415664 119494 415676
rect 137646 415664 137652 415676
rect 119488 415636 137652 415664
rect 119488 415624 119494 415636
rect 137646 415624 137652 415636
rect 137704 415624 137710 415676
rect 148318 415624 148324 415676
rect 148376 415664 148382 415676
rect 165706 415664 165712 415676
rect 148376 415636 165712 415664
rect 148376 415624 148382 415636
rect 165706 415624 165712 415636
rect 165764 415624 165770 415676
rect 175458 415624 175464 415676
rect 175516 415664 175522 415676
rect 193674 415664 193680 415676
rect 175516 415636 193680 415664
rect 175516 415624 175522 415636
rect 193674 415624 193680 415636
rect 193732 415624 193738 415676
rect 203518 415624 203524 415676
rect 203576 415664 203582 415676
rect 221366 415664 221372 415676
rect 203576 415636 221372 415664
rect 203576 415624 203582 415636
rect 221366 415624 221372 415636
rect 221424 415624 221430 415676
rect 408034 415624 408040 415676
rect 408092 415664 408098 415676
rect 428642 415664 428648 415676
rect 408092 415636 428648 415664
rect 408092 415624 408098 415636
rect 428642 415624 428648 415636
rect 428700 415624 428706 415676
rect 492030 415624 492036 415676
rect 492088 415664 492094 415676
rect 512730 415664 512736 415676
rect 492088 415636 512736 415664
rect 492088 415624 492094 415636
rect 512730 415624 512736 415636
rect 512788 415624 512794 415676
rect 36998 415556 37004 415608
rect 37056 415596 37062 415608
rect 53650 415596 53656 415608
rect 37056 415568 53656 415596
rect 37056 415556 37062 415568
rect 53650 415556 53656 415568
rect 53708 415556 53714 415608
rect 64322 415556 64328 415608
rect 64380 415596 64386 415608
rect 81434 415596 81440 415608
rect 64380 415568 81440 415596
rect 64380 415556 64386 415568
rect 81434 415556 81440 415568
rect 81492 415556 81498 415608
rect 91462 415556 91468 415608
rect 91520 415596 91526 415608
rect 109678 415596 109684 415608
rect 91520 415568 109684 415596
rect 91520 415556 91526 415568
rect 109678 415556 109684 415568
rect 109736 415556 109742 415608
rect 127986 415556 127992 415608
rect 128044 415596 128050 415608
rect 148502 415596 148508 415608
rect 128044 415568 148508 415596
rect 128044 415556 128050 415568
rect 148502 415556 148508 415568
rect 148560 415556 148566 415608
rect 156322 415556 156328 415608
rect 156380 415596 156386 415608
rect 178678 415596 178684 415608
rect 156380 415568 178684 415596
rect 156380 415556 156386 415568
rect 178678 415556 178684 415568
rect 178736 415556 178742 415608
rect 232590 415556 232596 415608
rect 232648 415596 232654 415608
rect 249702 415596 249708 415608
rect 232648 415568 249708 415596
rect 232648 415556 232654 415568
rect 249702 415556 249708 415568
rect 249760 415556 249766 415608
rect 260190 415556 260196 415608
rect 260248 415596 260254 415608
rect 277670 415596 277676 415608
rect 260248 415568 277676 415596
rect 260248 415556 260254 415568
rect 277670 415556 277676 415568
rect 277728 415556 277734 415608
rect 287514 415556 287520 415608
rect 287572 415596 287578 415608
rect 305362 415596 305368 415608
rect 287572 415568 305368 415596
rect 287572 415556 287578 415568
rect 305362 415556 305368 415568
rect 305420 415556 305426 415608
rect 315482 415556 315488 415608
rect 315540 415596 315546 415608
rect 333698 415596 333704 415608
rect 315540 415568 333704 415596
rect 315540 415556 315546 415568
rect 333698 415556 333704 415568
rect 333756 415556 333762 415608
rect 345658 415556 345664 415608
rect 345716 415596 345722 415608
rect 361666 415596 361672 415608
rect 345716 415568 361672 415596
rect 345716 415556 345722 415568
rect 361666 415556 361672 415568
rect 361724 415556 361730 415608
rect 371510 415556 371516 415608
rect 371568 415596 371574 415608
rect 389358 415596 389364 415608
rect 371568 415568 389364 415596
rect 371568 415556 371574 415568
rect 389358 415556 389364 415568
rect 389416 415556 389422 415608
rect 399478 415556 399484 415608
rect 399536 415596 399542 415608
rect 417694 415596 417700 415608
rect 399536 415568 417700 415596
rect 399536 415556 399542 415568
rect 417694 415556 417700 415568
rect 417752 415556 417758 415608
rect 456150 415556 456156 415608
rect 456208 415596 456214 415608
rect 473354 415596 473360 415608
rect 456208 415568 473360 415596
rect 456208 415556 456214 415568
rect 473354 415556 473360 415568
rect 473412 415556 473418 415608
rect 483474 415556 483480 415608
rect 483532 415596 483538 415608
rect 501690 415596 501696 415608
rect 483532 415568 501696 415596
rect 483532 415556 483538 415568
rect 501690 415556 501696 415568
rect 501748 415556 501754 415608
rect 36906 415488 36912 415540
rect 36964 415528 36970 415540
rect 63310 415528 63316 415540
rect 36964 415500 63316 415528
rect 36964 415488 36970 415500
rect 63310 415488 63316 415500
rect 63368 415488 63374 415540
rect 66898 415488 66904 415540
rect 66956 415528 66962 415540
rect 91094 415528 91100 415540
rect 66956 415500 91100 415528
rect 66956 415488 66962 415500
rect 91094 415488 91100 415500
rect 91152 415488 91158 415540
rect 94498 415488 94504 415540
rect 94556 415528 94562 415540
rect 119338 415528 119344 415540
rect 94556 415500 119344 415528
rect 94556 415488 94562 415500
rect 119338 415488 119344 415500
rect 119396 415488 119402 415540
rect 120718 415488 120724 415540
rect 120776 415528 120782 415540
rect 147306 415528 147312 415540
rect 120776 415500 147312 415528
rect 120776 415488 120782 415500
rect 147306 415488 147312 415500
rect 147364 415488 147370 415540
rect 148410 415488 148416 415540
rect 148468 415528 148474 415540
rect 175366 415528 175372 415540
rect 148468 415500 175372 415528
rect 148468 415488 148474 415500
rect 175366 415488 175372 415500
rect 175424 415488 175430 415540
rect 177298 415488 177304 415540
rect 177356 415528 177362 415540
rect 203334 415528 203340 415540
rect 177356 415500 203340 415528
rect 177356 415488 177362 415500
rect 203334 415488 203340 415500
rect 203392 415488 203398 415540
rect 204898 415488 204904 415540
rect 204956 415528 204962 415540
rect 231026 415528 231032 415540
rect 204956 415500 231032 415528
rect 204956 415488 204962 415500
rect 231026 415488 231032 415500
rect 231084 415488 231090 415540
rect 232498 415488 232504 415540
rect 232556 415528 232562 415540
rect 259362 415528 259368 415540
rect 232556 415500 259368 415528
rect 232556 415488 232562 415500
rect 259362 415488 259368 415500
rect 259420 415488 259426 415540
rect 268010 415488 268016 415540
rect 268068 415528 268074 415540
rect 287698 415528 287704 415540
rect 268068 415500 287704 415528
rect 268068 415488 268074 415500
rect 287698 415488 287704 415500
rect 287756 415488 287762 415540
rect 296346 415488 296352 415540
rect 296404 415528 296410 415540
rect 316770 415528 316776 415540
rect 296404 415500 316776 415528
rect 296404 415488 296410 415500
rect 316770 415488 316776 415500
rect 316828 415488 316834 415540
rect 352006 415488 352012 415540
rect 352064 415528 352070 415540
rect 374638 415528 374644 415540
rect 352064 415500 374644 415528
rect 352064 415488 352070 415500
rect 374638 415488 374644 415500
rect 374696 415488 374702 415540
rect 428550 415488 428556 415540
rect 428608 415528 428614 415540
rect 445662 415528 445668 415540
rect 428608 415500 445668 415528
rect 428608 415488 428614 415500
rect 445662 415488 445668 415500
rect 445720 415488 445726 415540
rect 464338 415488 464344 415540
rect 464396 415528 464402 415540
rect 483658 415528 483664 415540
rect 464396 415500 483664 415528
rect 464396 415488 464402 415500
rect 483658 415488 483664 415500
rect 483716 415488 483722 415540
rect 511442 415488 511448 415540
rect 511500 415528 511506 415540
rect 529658 415528 529664 415540
rect 511500 415500 529664 415528
rect 511500 415488 511506 415500
rect 529658 415488 529664 415500
rect 529716 415488 529722 415540
rect 542998 415488 543004 415540
rect 543056 415528 543062 415540
rect 557534 415528 557540 415540
rect 543056 415500 557540 415528
rect 543056 415488 543062 415500
rect 557534 415488 557540 415500
rect 557592 415488 557598 415540
rect 212350 415420 212356 415472
rect 212408 415460 212414 415472
rect 232682 415460 232688 415472
rect 212408 415432 232688 415460
rect 212408 415420 212414 415432
rect 232682 415420 232688 415432
rect 232740 415420 232746 415472
rect 260098 415420 260104 415472
rect 260156 415460 260162 415472
rect 287330 415460 287336 415472
rect 260156 415432 287336 415460
rect 260156 415420 260162 415432
rect 287330 415420 287336 415432
rect 287388 415420 287394 415472
rect 289078 415420 289084 415472
rect 289136 415460 289142 415472
rect 315022 415460 315028 415472
rect 289136 415432 315028 415460
rect 289136 415420 289142 415432
rect 315022 415420 315028 415432
rect 315080 415420 315086 415472
rect 316678 415420 316684 415472
rect 316736 415460 316742 415472
rect 343358 415460 343364 415472
rect 316736 415432 343364 415460
rect 316736 415420 316742 415432
rect 343358 415420 343364 415432
rect 343416 415420 343422 415472
rect 344278 415420 344284 415472
rect 344336 415460 344342 415472
rect 371326 415460 371332 415472
rect 344336 415432 371332 415460
rect 344336 415420 344342 415432
rect 371326 415420 371332 415432
rect 371384 415420 371390 415472
rect 373258 415420 373264 415472
rect 373316 415460 373322 415472
rect 399018 415460 399024 415472
rect 373316 415432 399024 415460
rect 373316 415420 373322 415432
rect 399018 415420 399024 415432
rect 399076 415420 399082 415472
rect 400858 415420 400864 415472
rect 400916 415460 400922 415472
rect 427354 415460 427360 415472
rect 400916 415432 427360 415460
rect 400916 415420 400922 415432
rect 427354 415420 427360 415432
rect 427412 415420 427418 415472
rect 428458 415420 428464 415472
rect 428516 415460 428522 415472
rect 455322 415460 455328 415472
rect 428516 415432 455328 415460
rect 428516 415420 428522 415432
rect 455322 415420 455328 415432
rect 455380 415420 455386 415472
rect 456058 415420 456064 415472
rect 456116 415460 456122 415472
rect 483014 415460 483020 415472
rect 456116 415432 483020 415460
rect 456116 415420 456122 415432
rect 483014 415420 483020 415432
rect 483072 415420 483078 415472
rect 485038 415420 485044 415472
rect 485096 415460 485102 415472
rect 511350 415460 511356 415472
rect 485096 415432 511356 415460
rect 485096 415420 485102 415432
rect 511350 415420 511356 415432
rect 511408 415420 511414 415472
rect 512638 415420 512644 415472
rect 512696 415460 512702 415472
rect 539318 415460 539324 415472
rect 512696 415432 539324 415460
rect 512696 415420 512702 415432
rect 539318 415420 539324 415432
rect 539376 415420 539382 415472
rect 540238 415420 540244 415472
rect 540296 415460 540302 415472
rect 567194 415460 567200 415472
rect 540296 415432 567200 415460
rect 540296 415420 540302 415432
rect 567194 415420 567200 415432
rect 567252 415420 567258 415472
rect 37918 414672 37924 414724
rect 37976 414712 37982 414724
rect 545758 414712 545764 414724
rect 37976 414684 545764 414712
rect 37976 414672 37982 414684
rect 545758 414672 545764 414684
rect 545816 414672 545822 414724
rect 35618 412632 35624 412684
rect 35676 412672 35682 412684
rect 36814 412672 36820 412684
rect 35676 412644 36820 412672
rect 35676 412632 35682 412644
rect 36814 412632 36820 412644
rect 36872 412632 36878 412684
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 13078 409884 13084 409896
rect 3384 409856 13084 409884
rect 3384 409844 3390 409856
rect 13078 409844 13084 409856
rect 13136 409844 13142 409896
rect 259730 398488 259736 398540
rect 259788 398528 259794 398540
rect 260190 398528 260196 398540
rect 259788 398500 260196 398528
rect 259788 398488 259794 398500
rect 260190 398488 260196 398500
rect 260248 398488 260254 398540
rect 455690 398488 455696 398540
rect 455748 398528 455754 398540
rect 456150 398528 456156 398540
rect 455748 398500 456156 398528
rect 455748 398488 455754 398500
rect 456150 398488 456156 398500
rect 456208 398488 456214 398540
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 11698 397508 11704 397520
rect 3384 397480 11704 397508
rect 3384 397468 3390 397480
rect 11698 397468 11704 397480
rect 11756 397468 11762 397520
rect 148502 395292 148508 395344
rect 148560 395332 148566 395344
rect 155862 395332 155868 395344
rect 148560 395304 155868 395332
rect 148560 395292 148566 395304
rect 155862 395292 155868 395304
rect 155920 395292 155926 395344
rect 428642 395292 428648 395344
rect 428700 395332 428706 395344
rect 435726 395332 435732 395344
rect 428700 395304 435732 395332
rect 428700 395292 428706 395304
rect 435726 395292 435732 395304
rect 435784 395292 435790 395344
rect 287698 395088 287704 395140
rect 287756 395128 287762 395140
rect 295794 395128 295800 395140
rect 287756 395100 295800 395128
rect 287756 395088 287762 395100
rect 295794 395088 295800 395100
rect 295852 395088 295858 395140
rect 316770 395088 316776 395140
rect 316828 395128 316834 395140
rect 323670 395128 323676 395140
rect 316828 395100 323676 395128
rect 316828 395088 316834 395100
rect 323670 395088 323676 395100
rect 323728 395088 323734 395140
rect 232682 395020 232688 395072
rect 232740 395060 232746 395072
rect 239766 395060 239772 395072
rect 232740 395032 239772 395060
rect 232740 395020 232746 395032
rect 239766 395020 239772 395032
rect 239824 395020 239830 395072
rect 483658 395020 483664 395072
rect 483716 395060 483722 395072
rect 491662 395060 491668 395072
rect 483716 395032 491668 395060
rect 483716 395020 483722 395032
rect 491662 395020 491668 395032
rect 491720 395020 491726 395072
rect 512730 395020 512736 395072
rect 512788 395060 512794 395072
rect 519630 395060 519636 395072
rect 512788 395032 519636 395060
rect 512788 395020 512794 395032
rect 519630 395020 519636 395032
rect 519688 395020 519694 395072
rect 13722 394612 13728 394664
rect 13780 394652 13786 394664
rect 13780 394624 59952 394652
rect 13780 394612 13786 394624
rect 35618 394544 35624 394596
rect 35676 394584 35682 394596
rect 36998 394584 37004 394596
rect 35676 394556 37004 394584
rect 35676 394544 35682 394556
rect 36998 394544 37004 394556
rect 37056 394544 37062 394596
rect 42702 394544 42708 394596
rect 42760 394584 42766 394596
rect 42760 394556 45554 394584
rect 42760 394544 42766 394556
rect 45526 394448 45554 394556
rect 59924 394516 59952 394624
rect 63586 394612 63592 394664
rect 63644 394652 63650 394664
rect 64322 394652 64328 394664
rect 63644 394624 64328 394652
rect 63644 394612 63650 394624
rect 64322 394612 64328 394624
rect 64380 394612 64386 394664
rect 70302 394612 70308 394664
rect 70360 394652 70366 394664
rect 121454 394652 121460 394664
rect 70360 394624 121460 394652
rect 70360 394612 70366 394624
rect 121454 394612 121460 394624
rect 121512 394612 121518 394664
rect 126882 394612 126888 394664
rect 126940 394652 126946 394664
rect 178034 394652 178040 394664
rect 126940 394624 178040 394652
rect 126940 394612 126946 394624
rect 178034 394612 178040 394624
rect 178092 394612 178098 394664
rect 209682 394612 209688 394664
rect 209740 394652 209746 394664
rect 262214 394652 262220 394664
rect 209740 394624 262220 394652
rect 209740 394612 209746 394624
rect 262214 394612 262220 394624
rect 262272 394612 262278 394664
rect 266262 394612 266268 394664
rect 266320 394652 266326 394664
rect 317414 394652 317420 394664
rect 266320 394624 317420 394652
rect 266320 394612 266326 394624
rect 317414 394612 317420 394624
rect 317472 394612 317478 394664
rect 322842 394612 322848 394664
rect 322900 394652 322906 394664
rect 373994 394652 374000 394664
rect 322900 394624 374000 394652
rect 322900 394612 322906 394624
rect 373994 394612 374000 394624
rect 374052 394612 374058 394664
rect 405642 394612 405648 394664
rect 405700 394652 405706 394664
rect 458174 394652 458180 394664
rect 405700 394624 458180 394652
rect 405700 394612 405706 394624
rect 458174 394612 458180 394624
rect 458232 394612 458238 394664
rect 489822 394612 489828 394664
rect 489880 394652 489886 394664
rect 542354 394652 542360 394664
rect 489880 394624 542360 394652
rect 489880 394612 489886 394624
rect 542354 394612 542360 394624
rect 542412 394612 542418 394664
rect 93854 394584 93860 394596
rect 74506 394556 93860 394584
rect 66254 394516 66260 394528
rect 59924 394488 66260 394516
rect 66254 394476 66260 394488
rect 66312 394476 66318 394528
rect 74506 394448 74534 394556
rect 93854 394544 93860 394556
rect 93912 394544 93918 394596
rect 97902 394544 97908 394596
rect 97960 394584 97966 394596
rect 149054 394584 149060 394596
rect 97960 394556 149060 394584
rect 97960 394544 97966 394556
rect 149054 394544 149060 394556
rect 149112 394544 149118 394596
rect 182082 394544 182088 394596
rect 182140 394584 182146 394596
rect 233234 394584 233240 394596
rect 182140 394556 233240 394584
rect 182140 394544 182146 394556
rect 233234 394544 233240 394556
rect 233292 394544 233298 394596
rect 238662 394544 238668 394596
rect 238720 394584 238726 394596
rect 289814 394584 289820 394596
rect 238720 394556 289820 394584
rect 238720 394544 238726 394556
rect 289814 394544 289820 394556
rect 289872 394544 289878 394596
rect 293862 394544 293868 394596
rect 293920 394584 293926 394596
rect 293920 394556 335354 394584
rect 293920 394544 293926 394556
rect 154482 394476 154488 394528
rect 154540 394516 154546 394528
rect 205634 394516 205640 394528
rect 154540 394488 205640 394516
rect 154540 394476 154546 394488
rect 205634 394476 205640 394488
rect 205692 394476 205698 394528
rect 335326 394516 335354 394556
rect 343634 394544 343640 394596
rect 343692 394584 343698 394596
rect 345658 394584 345664 394596
rect 343692 394556 345664 394584
rect 343692 394544 343698 394556
rect 345658 394544 345664 394556
rect 345716 394544 345722 394596
rect 350442 394544 350448 394596
rect 350500 394584 350506 394596
rect 401594 394584 401600 394596
rect 350500 394556 401600 394584
rect 350500 394544 350506 394556
rect 401594 394544 401600 394556
rect 401652 394544 401658 394596
rect 427722 394544 427728 394596
rect 427780 394584 427786 394596
rect 428550 394584 428556 394596
rect 427780 394556 428556 394584
rect 427780 394544 427786 394556
rect 428550 394544 428556 394556
rect 428608 394544 428614 394596
rect 462222 394544 462228 394596
rect 462280 394584 462286 394596
rect 513374 394584 513380 394596
rect 462280 394556 513380 394584
rect 462280 394544 462286 394556
rect 513374 394544 513380 394556
rect 513432 394544 513438 394596
rect 518802 394544 518808 394596
rect 518860 394584 518866 394596
rect 569954 394584 569960 394596
rect 518860 394556 569960 394584
rect 518860 394544 518866 394556
rect 569954 394544 569960 394556
rect 570012 394544 570018 394596
rect 345014 394516 345020 394528
rect 335326 394488 345020 394516
rect 345014 394476 345020 394488
rect 345072 394476 345078 394528
rect 378042 394476 378048 394528
rect 378100 394516 378106 394528
rect 429194 394516 429200 394528
rect 378100 394488 429200 394516
rect 378100 394476 378106 394488
rect 429194 394476 429200 394488
rect 429252 394476 429258 394528
rect 434622 394476 434628 394528
rect 434680 394516 434686 394528
rect 485774 394516 485780 394528
rect 434680 394488 485780 394516
rect 434680 394476 434686 394488
rect 485774 394476 485780 394488
rect 485832 394476 485838 394528
rect 45526 394420 74534 394448
rect 231578 393252 231584 393304
rect 231636 393292 231642 393304
rect 232590 393292 232596 393304
rect 231636 393264 232596 393292
rect 231636 393252 231642 393264
rect 232590 393252 232596 393264
rect 232648 393252 232654 393304
rect 25682 391892 25688 391944
rect 25740 391932 25746 391944
rect 36906 391932 36912 391944
rect 25740 391904 36912 391932
rect 25740 391892 25746 391904
rect 36906 391892 36912 391904
rect 36964 391892 36970 391944
rect 178678 391892 178684 391944
rect 178736 391932 178742 391944
rect 184014 391932 184020 391944
rect 178736 391904 184020 391932
rect 178736 391892 178742 391904
rect 184014 391892 184020 391904
rect 184072 391892 184078 391944
rect 374638 391892 374644 391944
rect 374696 391932 374702 391944
rect 379698 391932 379704 391944
rect 374696 391904 379704 391932
rect 374696 391892 374702 391904
rect 379698 391892 379704 391904
rect 379756 391892 379762 391944
rect 539318 391892 539324 391944
rect 539376 391932 539382 391944
rect 542998 391932 543004 391944
rect 539376 391904 543004 391932
rect 539376 391892 539382 391904
rect 542998 391892 543004 391904
rect 543056 391892 543062 391944
rect 15194 391824 15200 391876
rect 15252 391864 15258 391876
rect 43990 391864 43996 391876
rect 15252 391836 43996 391864
rect 15252 391824 15258 391836
rect 43990 391824 43996 391836
rect 44048 391824 44054 391876
rect 69658 391824 69664 391876
rect 69716 391864 69722 391876
rect 567194 391864 567200 391876
rect 69716 391836 567200 391864
rect 69716 391824 69722 391836
rect 567194 391824 567200 391836
rect 567252 391824 567258 391876
rect 53650 391756 53656 391808
rect 53708 391796 53714 391808
rect 66898 391796 66904 391808
rect 53708 391768 66904 391796
rect 53708 391756 53714 391768
rect 66898 391756 66904 391768
rect 66956 391756 66962 391808
rect 71866 391756 71872 391808
rect 71924 391796 71930 391808
rect 100018 391796 100024 391808
rect 71924 391768 100024 391796
rect 71924 391756 71930 391768
rect 100018 391756 100024 391768
rect 100076 391756 100082 391808
rect 127986 391796 127992 391808
rect 103486 391768 127992 391796
rect 42886 391688 42892 391740
rect 42944 391728 42950 391740
rect 71958 391728 71964 391740
rect 42944 391700 71964 391728
rect 42944 391688 42950 391700
rect 71958 391688 71964 391700
rect 72016 391688 72022 391740
rect 81986 391688 81992 391740
rect 82044 391728 82050 391740
rect 94498 391728 94504 391740
rect 82044 391700 94504 391728
rect 82044 391688 82050 391700
rect 94498 391688 94504 391700
rect 94556 391688 94562 391740
rect 99466 391688 99472 391740
rect 99524 391728 99530 391740
rect 103486 391728 103514 391768
rect 127986 391756 127992 391768
rect 128044 391756 128050 391808
rect 137646 391756 137652 391808
rect 137704 391796 137710 391808
rect 148410 391796 148416 391808
rect 137704 391768 148416 391796
rect 137704 391756 137710 391768
rect 148410 391756 148416 391768
rect 148468 391756 148474 391808
rect 165982 391756 165988 391808
rect 166040 391796 166046 391808
rect 177298 391796 177304 391808
rect 166040 391768 177304 391796
rect 166040 391756 166046 391768
rect 177298 391756 177304 391768
rect 177356 391756 177362 391808
rect 183646 391756 183652 391808
rect 183704 391796 183710 391808
rect 211706 391796 211712 391808
rect 183704 391768 211712 391796
rect 183704 391756 183710 391768
rect 211706 391756 211712 391768
rect 211764 391756 211770 391808
rect 221918 391756 221924 391808
rect 221976 391796 221982 391808
rect 232498 391796 232504 391808
rect 221976 391768 232504 391796
rect 221976 391756 221982 391768
rect 232498 391756 232504 391768
rect 232556 391756 232562 391808
rect 238846 391756 238852 391808
rect 238904 391796 238910 391808
rect 268010 391796 268016 391808
rect 238904 391768 268016 391796
rect 238904 391756 238910 391768
rect 268010 391756 268016 391768
rect 268068 391756 268074 391808
rect 277670 391756 277676 391808
rect 277728 391796 277734 391808
rect 289078 391796 289084 391808
rect 277728 391768 289084 391796
rect 277728 391756 277734 391768
rect 289078 391756 289084 391768
rect 289136 391756 289142 391808
rect 306006 391756 306012 391808
rect 306064 391796 306070 391808
rect 316678 391796 316684 391808
rect 306064 391768 316684 391796
rect 306064 391756 306070 391768
rect 316678 391756 316684 391768
rect 316736 391756 316742 391808
rect 323026 391756 323032 391808
rect 323084 391796 323090 391808
rect 352006 391796 352012 391808
rect 323084 391768 352012 391796
rect 323084 391756 323090 391768
rect 352006 391756 352012 391768
rect 352064 391756 352070 391808
rect 361666 391756 361672 391808
rect 361724 391796 361730 391808
rect 373258 391796 373264 391808
rect 361724 391768 373264 391796
rect 361724 391756 361730 391768
rect 373258 391756 373264 391768
rect 373316 391756 373322 391808
rect 379606 391756 379612 391808
rect 379664 391796 379670 391808
rect 408034 391796 408040 391808
rect 379664 391768 408040 391796
rect 379664 391756 379670 391768
rect 408034 391756 408040 391768
rect 408092 391756 408098 391808
rect 417694 391756 417700 391808
rect 417752 391796 417758 391808
rect 428458 391796 428464 391808
rect 417752 391768 428464 391796
rect 417752 391756 417758 391768
rect 428458 391756 428464 391768
rect 428516 391756 428522 391808
rect 434806 391756 434812 391808
rect 434864 391796 434870 391808
rect 463786 391796 463792 391808
rect 434864 391768 463792 391796
rect 434864 391756 434870 391768
rect 463786 391756 463792 391768
rect 463844 391756 463850 391808
rect 473998 391756 474004 391808
rect 474056 391796 474062 391808
rect 485038 391796 485044 391808
rect 474056 391768 485044 391796
rect 474056 391756 474062 391768
rect 485038 391756 485044 391768
rect 485096 391756 485102 391808
rect 501690 391756 501696 391808
rect 501748 391796 501754 391808
rect 512638 391796 512644 391808
rect 501748 391768 512644 391796
rect 501748 391756 501754 391768
rect 512638 391756 512644 391768
rect 512696 391756 512702 391808
rect 518986 391756 518992 391808
rect 519044 391796 519050 391808
rect 547874 391796 547880 391808
rect 519044 391768 547880 391796
rect 519044 391756 519050 391768
rect 547874 391756 547880 391768
rect 547932 391756 547938 391808
rect 99524 391700 103514 391728
rect 99524 391688 99530 391700
rect 109678 391688 109684 391740
rect 109736 391728 109742 391740
rect 120718 391728 120724 391740
rect 109736 391700 120724 391728
rect 109736 391688 109742 391700
rect 120718 391688 120724 391700
rect 120776 391688 120782 391740
rect 193674 391688 193680 391740
rect 193732 391728 193738 391740
rect 204898 391728 204904 391740
rect 193732 391700 204904 391728
rect 193732 391688 193738 391700
rect 204898 391688 204904 391700
rect 204956 391688 204962 391740
rect 249702 391688 249708 391740
rect 249760 391728 249766 391740
rect 260098 391728 260104 391740
rect 249760 391700 260104 391728
rect 249760 391688 249766 391700
rect 260098 391688 260104 391700
rect 260156 391688 260162 391740
rect 333698 391688 333704 391740
rect 333756 391728 333762 391740
rect 344278 391728 344284 391740
rect 333756 391700 344284 391728
rect 333756 391688 333762 391700
rect 344278 391688 344284 391700
rect 344336 391688 344342 391740
rect 390002 391688 390008 391740
rect 390060 391728 390066 391740
rect 400858 391728 400864 391740
rect 390060 391700 400864 391728
rect 390060 391688 390066 391700
rect 400858 391688 400864 391700
rect 400916 391688 400922 391740
rect 445662 391688 445668 391740
rect 445720 391728 445726 391740
rect 456058 391728 456064 391740
rect 445720 391700 456064 391728
rect 445720 391688 445726 391700
rect 456058 391688 456064 391700
rect 456116 391688 456122 391740
rect 529658 391688 529664 391740
rect 529716 391728 529722 391740
rect 540238 391728 540244 391740
rect 529716 391700 540244 391728
rect 529716 391688 529722 391700
rect 540238 391688 540244 391700
rect 540296 391688 540302 391740
rect 36722 391620 36728 391672
rect 36780 391660 36786 391672
rect 557534 391660 557540 391672
rect 36780 391632 557540 391660
rect 36780 391620 36786 391632
rect 557534 391620 557540 391632
rect 557592 391620 557598 391672
rect 16022 389784 16028 389836
rect 16080 389824 16086 389836
rect 547874 389824 547880 389836
rect 16080 389796 547880 389824
rect 16080 389784 16086 389796
rect 547874 389784 547880 389796
rect 547932 389784 547938 389836
rect 25682 389376 25688 389428
rect 25740 389416 25746 389428
rect 71038 389416 71044 389428
rect 25740 389388 71044 389416
rect 25740 389376 25746 389388
rect 71038 389376 71044 389388
rect 71096 389376 71102 389428
rect 212350 389376 212356 389428
rect 212408 389416 212414 389428
rect 232682 389416 232688 389428
rect 212408 389388 232688 389416
rect 212408 389376 212414 389388
rect 232682 389376 232688 389388
rect 232740 389376 232746 389428
rect 296346 389376 296352 389428
rect 296404 389416 296410 389428
rect 316770 389416 316776 389428
rect 296404 389388 316776 389416
rect 296404 389376 296410 389388
rect 316770 389376 316776 389388
rect 316828 389376 316834 389428
rect 408034 389376 408040 389428
rect 408092 389416 408098 389428
rect 428642 389416 428648 389428
rect 408092 389388 428648 389416
rect 408092 389376 408098 389388
rect 428642 389376 428648 389388
rect 428700 389376 428706 389428
rect 492030 389376 492036 389428
rect 492088 389416 492094 389428
rect 512730 389416 512736 389428
rect 492088 389388 512736 389416
rect 492088 389376 492094 389388
rect 512730 389376 512736 389388
rect 512788 389376 512794 389428
rect 36998 389308 37004 389360
rect 37056 389348 37062 389360
rect 53650 389348 53656 389360
rect 37056 389320 53656 389348
rect 37056 389308 37062 389320
rect 53650 389308 53656 389320
rect 53708 389308 53714 389360
rect 148410 389308 148416 389360
rect 148468 389348 148474 389360
rect 165706 389348 165712 389360
rect 148468 389320 165712 389348
rect 148468 389308 148474 389320
rect 165706 389308 165712 389320
rect 165764 389308 165770 389360
rect 175458 389308 175464 389360
rect 175516 389348 175522 389360
rect 193674 389348 193680 389360
rect 175516 389320 193680 389348
rect 175516 389308 175522 389320
rect 193674 389308 193680 389320
rect 193732 389308 193738 389360
rect 203518 389308 203524 389360
rect 203576 389348 203582 389360
rect 221366 389348 221372 389360
rect 203576 389320 221372 389348
rect 203576 389308 203582 389320
rect 221366 389308 221372 389320
rect 221424 389308 221430 389360
rect 260098 389308 260104 389360
rect 260156 389348 260162 389360
rect 277670 389348 277676 389360
rect 260156 389320 277676 389348
rect 260156 389308 260162 389320
rect 277670 389308 277676 389320
rect 277728 389308 277734 389360
rect 287514 389308 287520 389360
rect 287572 389348 287578 389360
rect 305362 389348 305368 389360
rect 287572 389320 305368 389348
rect 287572 389308 287578 389320
rect 305362 389308 305368 389320
rect 305420 389308 305426 389360
rect 345658 389308 345664 389360
rect 345716 389348 345722 389360
rect 361666 389348 361672 389360
rect 345716 389320 361672 389348
rect 345716 389308 345722 389320
rect 361666 389308 361672 389320
rect 361724 389308 361730 389360
rect 371510 389308 371516 389360
rect 371568 389348 371574 389360
rect 389358 389348 389364 389360
rect 371568 389320 389364 389348
rect 371568 389308 371574 389320
rect 389358 389308 389364 389320
rect 389416 389308 389422 389360
rect 399478 389308 399484 389360
rect 399536 389348 399542 389360
rect 417694 389348 417700 389360
rect 399536 389320 417700 389348
rect 399536 389308 399542 389320
rect 417694 389308 417700 389320
rect 417752 389308 417758 389360
rect 456150 389308 456156 389360
rect 456208 389348 456214 389360
rect 473354 389348 473360 389360
rect 456208 389320 473360 389348
rect 456208 389308 456214 389320
rect 473354 389308 473360 389320
rect 473412 389308 473418 389360
rect 483474 389308 483480 389360
rect 483532 389348 483538 389360
rect 501690 389348 501696 389360
rect 483532 389320 501696 389348
rect 483532 389308 483538 389320
rect 501690 389308 501696 389320
rect 501748 389308 501754 389360
rect 36906 389240 36912 389292
rect 36964 389280 36970 389292
rect 63310 389280 63316 389292
rect 36964 389252 63316 389280
rect 36964 389240 36970 389252
rect 63310 389240 63316 389252
rect 63368 389240 63374 389292
rect 64322 389240 64328 389292
rect 64380 389280 64386 389292
rect 81434 389280 81440 389292
rect 64380 389252 81440 389280
rect 64380 389240 64386 389252
rect 81434 389240 81440 389252
rect 81492 389240 81498 389292
rect 91462 389240 91468 389292
rect 91520 389280 91526 389292
rect 109678 389280 109684 389292
rect 91520 389252 109684 389280
rect 91520 389240 91526 389252
rect 109678 389240 109684 389252
rect 109736 389240 109742 389292
rect 119430 389240 119436 389292
rect 119488 389280 119494 389292
rect 137646 389280 137652 389292
rect 119488 389252 137652 389280
rect 119488 389240 119494 389252
rect 137646 389240 137652 389252
rect 137704 389240 137710 389292
rect 156322 389240 156328 389292
rect 156380 389280 156386 389292
rect 178678 389280 178684 389292
rect 156380 389252 178684 389280
rect 156380 389240 156386 389252
rect 178678 389240 178684 389252
rect 178736 389240 178742 389292
rect 232590 389240 232596 389292
rect 232648 389280 232654 389292
rect 249702 389280 249708 389292
rect 232648 389252 249708 389280
rect 232648 389240 232654 389252
rect 249702 389240 249708 389252
rect 249760 389240 249766 389292
rect 268010 389240 268016 389292
rect 268068 389280 268074 389292
rect 287698 389280 287704 389292
rect 268068 389252 287704 389280
rect 268068 389240 268074 389252
rect 287698 389240 287704 389252
rect 287756 389240 287762 389292
rect 315482 389240 315488 389292
rect 315540 389280 315546 389292
rect 333698 389280 333704 389292
rect 315540 389252 333704 389280
rect 315540 389240 315546 389252
rect 333698 389240 333704 389252
rect 333756 389240 333762 389292
rect 352006 389240 352012 389292
rect 352064 389280 352070 389292
rect 374638 389280 374644 389292
rect 352064 389252 374644 389280
rect 352064 389240 352070 389252
rect 374638 389240 374644 389252
rect 374696 389240 374702 389292
rect 428550 389240 428556 389292
rect 428608 389280 428614 389292
rect 445662 389280 445668 389292
rect 428608 389252 445668 389280
rect 428608 389240 428614 389252
rect 445662 389240 445668 389252
rect 445720 389240 445726 389292
rect 464338 389240 464344 389292
rect 464396 389280 464402 389292
rect 483658 389280 483664 389292
rect 464396 389252 483664 389280
rect 464396 389240 464402 389252
rect 483658 389240 483664 389252
rect 483716 389240 483722 389292
rect 511442 389240 511448 389292
rect 511500 389280 511506 389292
rect 529658 389280 529664 389292
rect 511500 389252 529664 389280
rect 511500 389240 511506 389252
rect 529658 389240 529664 389252
rect 529716 389240 529722 389292
rect 542998 389240 543004 389292
rect 543056 389280 543062 389292
rect 557534 389280 557540 389292
rect 543056 389252 557540 389280
rect 543056 389240 543062 389252
rect 557534 389240 557540 389252
rect 557592 389240 557598 389292
rect 69658 389172 69664 389224
rect 69716 389212 69722 389224
rect 91094 389212 91100 389224
rect 69716 389184 91100 389212
rect 69716 389172 69722 389184
rect 91094 389172 91100 389184
rect 91152 389172 91158 389224
rect 94498 389172 94504 389224
rect 94556 389212 94562 389224
rect 119338 389212 119344 389224
rect 94556 389184 119344 389212
rect 94556 389172 94562 389184
rect 119338 389172 119344 389184
rect 119396 389172 119402 389224
rect 120718 389172 120724 389224
rect 120776 389212 120782 389224
rect 147306 389212 147312 389224
rect 120776 389184 147312 389212
rect 120776 389172 120782 389184
rect 147306 389172 147312 389184
rect 147364 389172 147370 389224
rect 148318 389172 148324 389224
rect 148376 389212 148382 389224
rect 175366 389212 175372 389224
rect 148376 389184 175372 389212
rect 148376 389172 148382 389184
rect 175366 389172 175372 389184
rect 175424 389172 175430 389224
rect 177298 389172 177304 389224
rect 177356 389212 177362 389224
rect 203334 389212 203340 389224
rect 177356 389184 203340 389212
rect 177356 389172 177362 389184
rect 203334 389172 203340 389184
rect 203392 389172 203398 389224
rect 204898 389172 204904 389224
rect 204956 389212 204962 389224
rect 231026 389212 231032 389224
rect 204956 389184 231032 389212
rect 204956 389172 204962 389184
rect 231026 389172 231032 389184
rect 231084 389172 231090 389224
rect 232498 389172 232504 389224
rect 232556 389212 232562 389224
rect 259362 389212 259368 389224
rect 232556 389184 259368 389212
rect 232556 389172 232562 389184
rect 259362 389172 259368 389184
rect 259420 389172 259426 389224
rect 260190 389172 260196 389224
rect 260248 389212 260254 389224
rect 287330 389212 287336 389224
rect 260248 389184 287336 389212
rect 260248 389172 260254 389184
rect 287330 389172 287336 389184
rect 287388 389172 287394 389224
rect 289078 389172 289084 389224
rect 289136 389212 289142 389224
rect 315022 389212 315028 389224
rect 289136 389184 315028 389212
rect 289136 389172 289142 389184
rect 315022 389172 315028 389184
rect 315080 389172 315086 389224
rect 316678 389172 316684 389224
rect 316736 389212 316742 389224
rect 343358 389212 343364 389224
rect 316736 389184 343364 389212
rect 316736 389172 316742 389184
rect 343358 389172 343364 389184
rect 343416 389172 343422 389224
rect 344278 389172 344284 389224
rect 344336 389212 344342 389224
rect 371326 389212 371332 389224
rect 344336 389184 371332 389212
rect 344336 389172 344342 389184
rect 371326 389172 371332 389184
rect 371384 389172 371390 389224
rect 373258 389172 373264 389224
rect 373316 389212 373322 389224
rect 399018 389212 399024 389224
rect 373316 389184 399024 389212
rect 373316 389172 373322 389184
rect 399018 389172 399024 389184
rect 399076 389172 399082 389224
rect 400858 389172 400864 389224
rect 400916 389212 400922 389224
rect 427354 389212 427360 389224
rect 400916 389184 427360 389212
rect 400916 389172 400922 389184
rect 427354 389172 427360 389184
rect 427412 389172 427418 389224
rect 428458 389172 428464 389224
rect 428516 389212 428522 389224
rect 455322 389212 455328 389224
rect 428516 389184 455328 389212
rect 428516 389172 428522 389184
rect 455322 389172 455328 389184
rect 455380 389172 455386 389224
rect 456058 389172 456064 389224
rect 456116 389212 456122 389224
rect 483014 389212 483020 389224
rect 456116 389184 483020 389212
rect 456116 389172 456122 389184
rect 483014 389172 483020 389184
rect 483072 389172 483078 389224
rect 485038 389172 485044 389224
rect 485096 389212 485102 389224
rect 511350 389212 511356 389224
rect 485096 389184 511356 389212
rect 485096 389172 485102 389184
rect 511350 389172 511356 389184
rect 511408 389172 511414 389224
rect 512638 389172 512644 389224
rect 512696 389212 512702 389224
rect 539318 389212 539324 389224
rect 512696 389184 539324 389212
rect 512696 389172 512702 389184
rect 539318 389172 539324 389184
rect 539376 389172 539382 389224
rect 540238 389172 540244 389224
rect 540296 389212 540302 389224
rect 567194 389212 567200 389224
rect 540296 389184 567200 389212
rect 540296 389172 540302 389184
rect 567194 389172 567200 389184
rect 567252 389172 567258 389224
rect 37918 387064 37924 387116
rect 37976 387104 37982 387116
rect 545758 387104 545764 387116
rect 37976 387076 545764 387104
rect 37976 387064 37982 387076
rect 545758 387064 545764 387076
rect 545816 387064 545822 387116
rect 35618 386384 35624 386436
rect 35676 386424 35682 386436
rect 36722 386424 36728 386436
rect 35676 386396 36728 386424
rect 35676 386384 35682 386396
rect 36722 386384 36728 386396
rect 36780 386384 36786 386436
rect 63586 370540 63592 370592
rect 63644 370580 63650 370592
rect 64322 370580 64328 370592
rect 63644 370552 64328 370580
rect 63644 370540 63650 370552
rect 64322 370540 64328 370552
rect 64380 370540 64386 370592
rect 147674 370540 147680 370592
rect 147732 370580 147738 370592
rect 148410 370580 148416 370592
rect 147732 370552 148416 370580
rect 147732 370540 147738 370552
rect 148410 370540 148416 370552
rect 148468 370540 148474 370592
rect 455690 370540 455696 370592
rect 455748 370580 455754 370592
rect 456150 370580 456156 370592
rect 455748 370552 456156 370580
rect 455748 370540 455754 370552
rect 456150 370540 456156 370552
rect 456208 370540 456214 370592
rect 232682 369248 232688 369300
rect 232740 369288 232746 369300
rect 239766 369288 239772 369300
rect 232740 369260 239772 369288
rect 232740 369248 232746 369260
rect 239766 369248 239772 369260
rect 239824 369248 239830 369300
rect 428642 369112 428648 369164
rect 428700 369152 428706 369164
rect 435726 369152 435732 369164
rect 428700 369124 435732 369152
rect 428700 369112 428706 369124
rect 435726 369112 435732 369124
rect 435784 369112 435790 369164
rect 287698 368840 287704 368892
rect 287756 368880 287762 368892
rect 295702 368880 295708 368892
rect 287756 368852 295708 368880
rect 287756 368840 287762 368852
rect 295702 368840 295708 368852
rect 295760 368840 295766 368892
rect 316770 368840 316776 368892
rect 316828 368880 316834 368892
rect 323670 368880 323676 368892
rect 316828 368852 323676 368880
rect 316828 368840 316834 368852
rect 323670 368840 323676 368852
rect 323728 368840 323734 368892
rect 483658 368840 483664 368892
rect 483716 368880 483722 368892
rect 491662 368880 491668 368892
rect 483716 368852 491668 368880
rect 483716 368840 483722 368852
rect 491662 368840 491668 368852
rect 491720 368840 491726 368892
rect 512730 368704 512736 368756
rect 512788 368744 512794 368756
rect 519630 368744 519636 368756
rect 512788 368716 519636 368744
rect 512788 368704 512794 368716
rect 519630 368704 519636 368716
rect 519688 368704 519694 368756
rect 13722 368432 13728 368484
rect 13780 368472 13786 368484
rect 66254 368472 66260 368484
rect 13780 368444 66260 368472
rect 13780 368432 13786 368444
rect 66254 368432 66260 368444
rect 66312 368432 66318 368484
rect 70302 368432 70308 368484
rect 70360 368472 70366 368484
rect 121454 368472 121460 368484
rect 70360 368444 121460 368472
rect 70360 368432 70366 368444
rect 121454 368432 121460 368444
rect 121512 368432 121518 368484
rect 126882 368432 126888 368484
rect 126940 368472 126946 368484
rect 178034 368472 178040 368484
rect 126940 368444 178040 368472
rect 126940 368432 126946 368444
rect 178034 368432 178040 368444
rect 178092 368432 178098 368484
rect 209682 368432 209688 368484
rect 209740 368472 209746 368484
rect 260742 368472 260748 368484
rect 209740 368444 260748 368472
rect 209740 368432 209746 368444
rect 260742 368432 260748 368444
rect 260800 368432 260806 368484
rect 266262 368432 266268 368484
rect 266320 368472 266326 368484
rect 317414 368472 317420 368484
rect 266320 368444 317420 368472
rect 266320 368432 266326 368444
rect 317414 368432 317420 368444
rect 317472 368432 317478 368484
rect 322842 368432 322848 368484
rect 322900 368472 322906 368484
rect 373994 368472 374000 368484
rect 322900 368444 374000 368472
rect 322900 368432 322906 368444
rect 373994 368432 374000 368444
rect 374052 368432 374058 368484
rect 405642 368432 405648 368484
rect 405700 368472 405706 368484
rect 458174 368472 458180 368484
rect 405700 368444 458180 368472
rect 405700 368432 405706 368444
rect 458174 368432 458180 368444
rect 458232 368432 458238 368484
rect 489822 368432 489828 368484
rect 489880 368472 489886 368484
rect 540882 368472 540888 368484
rect 489880 368444 540888 368472
rect 489880 368432 489886 368444
rect 540882 368432 540888 368444
rect 540940 368432 540946 368484
rect 42702 368364 42708 368416
rect 42760 368404 42766 368416
rect 93854 368404 93860 368416
rect 42760 368376 93860 368404
rect 42760 368364 42766 368376
rect 93854 368364 93860 368376
rect 93912 368364 93918 368416
rect 97902 368364 97908 368416
rect 97960 368404 97966 368416
rect 149054 368404 149060 368416
rect 97960 368376 149060 368404
rect 97960 368364 97966 368376
rect 149054 368364 149060 368376
rect 149112 368364 149118 368416
rect 182082 368364 182088 368416
rect 182140 368404 182146 368416
rect 233234 368404 233240 368416
rect 182140 368376 233240 368404
rect 182140 368364 182146 368376
rect 233234 368364 233240 368376
rect 233292 368364 233298 368416
rect 238662 368364 238668 368416
rect 238720 368404 238726 368416
rect 289814 368404 289820 368416
rect 238720 368376 289820 368404
rect 238720 368364 238726 368376
rect 289814 368364 289820 368376
rect 289872 368364 289878 368416
rect 293862 368364 293868 368416
rect 293920 368404 293926 368416
rect 345014 368404 345020 368416
rect 293920 368376 345020 368404
rect 293920 368364 293926 368376
rect 345014 368364 345020 368376
rect 345072 368364 345078 368416
rect 378042 368364 378048 368416
rect 378100 368404 378106 368416
rect 429194 368404 429200 368416
rect 378100 368376 429200 368404
rect 378100 368364 378106 368376
rect 429194 368364 429200 368376
rect 429252 368364 429258 368416
rect 462222 368364 462228 368416
rect 462280 368404 462286 368416
rect 513374 368404 513380 368416
rect 462280 368376 513380 368404
rect 462280 368364 462286 368376
rect 513374 368364 513380 368376
rect 513432 368364 513438 368416
rect 518802 368364 518808 368416
rect 518860 368404 518866 368416
rect 569954 368404 569960 368416
rect 518860 368376 569960 368404
rect 518860 368364 518866 368376
rect 569954 368364 569960 368376
rect 570012 368364 570018 368416
rect 154482 368296 154488 368348
rect 154540 368336 154546 368348
rect 205634 368336 205640 368348
rect 154540 368308 205640 368336
rect 154540 368296 154546 368308
rect 205634 368296 205640 368308
rect 205692 368296 205698 368348
rect 231670 368296 231676 368348
rect 231728 368336 231734 368348
rect 232590 368336 232596 368348
rect 231728 368308 232596 368336
rect 231728 368296 231734 368308
rect 232590 368296 232596 368308
rect 232648 368296 232654 368348
rect 350442 368296 350448 368348
rect 350500 368336 350506 368348
rect 401594 368336 401600 368348
rect 350500 368308 401600 368336
rect 350500 368296 350506 368308
rect 401594 368296 401600 368308
rect 401652 368296 401658 368348
rect 427722 368296 427728 368348
rect 427780 368336 427786 368348
rect 428550 368336 428556 368348
rect 427780 368308 428556 368336
rect 427780 368296 427786 368308
rect 428550 368296 428556 368308
rect 428608 368296 428614 368348
rect 434622 368296 434628 368348
rect 434680 368336 434686 368348
rect 485774 368336 485780 368348
rect 434680 368308 485780 368336
rect 434680 368296 434686 368308
rect 485774 368296 485780 368308
rect 485832 368296 485838 368348
rect 35618 367004 35624 367056
rect 35676 367044 35682 367056
rect 36998 367044 37004 367056
rect 35676 367016 37004 367044
rect 35676 367004 35682 367016
rect 36998 367004 37004 367016
rect 37056 367004 37062 367056
rect 343542 367004 343548 367056
rect 343600 367044 343606 367056
rect 345658 367044 345664 367056
rect 343600 367016 345664 367044
rect 343600 367004 343606 367016
rect 345658 367004 345664 367016
rect 345716 367004 345722 367056
rect 25682 365644 25688 365696
rect 25740 365684 25746 365696
rect 36906 365684 36912 365696
rect 25740 365656 36912 365684
rect 25740 365644 25746 365656
rect 36906 365644 36912 365656
rect 36964 365644 36970 365696
rect 42886 365644 42892 365696
rect 42944 365684 42950 365696
rect 72050 365684 72056 365696
rect 42944 365656 45554 365684
rect 42944 365644 42950 365656
rect 15194 365576 15200 365628
rect 15252 365616 15258 365628
rect 43990 365616 43996 365628
rect 15252 365588 43996 365616
rect 15252 365576 15258 365588
rect 43990 365576 43996 365588
rect 44048 365576 44054 365628
rect 45526 365616 45554 365656
rect 64846 365656 72056 365684
rect 64846 365616 64874 365656
rect 72050 365644 72056 365656
rect 72108 365644 72114 365696
rect 99466 365644 99472 365696
rect 99524 365684 99530 365696
rect 99524 365656 103514 365684
rect 99524 365644 99530 365656
rect 45526 365588 64874 365616
rect 71866 365576 71872 365628
rect 71924 365616 71930 365628
rect 100018 365616 100024 365628
rect 71924 365588 100024 365616
rect 71924 365576 71930 365588
rect 100018 365576 100024 365588
rect 100076 365576 100082 365628
rect 103486 365616 103514 365656
rect 127066 365644 127072 365696
rect 127124 365684 127130 365696
rect 127124 365656 132494 365684
rect 127124 365644 127130 365656
rect 127986 365616 127992 365628
rect 103486 365588 127992 365616
rect 127986 365576 127992 365588
rect 128044 365576 128050 365628
rect 132466 365616 132494 365656
rect 183646 365644 183652 365696
rect 183704 365684 183710 365696
rect 183704 365656 190454 365684
rect 183704 365644 183710 365656
rect 156046 365616 156052 365628
rect 132466 365588 156052 365616
rect 156046 365576 156052 365588
rect 156104 365576 156110 365628
rect 165982 365576 165988 365628
rect 166040 365616 166046 365628
rect 177298 365616 177304 365628
rect 166040 365588 177304 365616
rect 166040 365576 166046 365588
rect 177298 365576 177304 365588
rect 177356 365576 177362 365628
rect 178678 365576 178684 365628
rect 178736 365616 178742 365628
rect 184014 365616 184020 365628
rect 178736 365588 184020 365616
rect 178736 365576 178742 365588
rect 184014 365576 184020 365588
rect 184072 365576 184078 365628
rect 190426 365616 190454 365656
rect 374638 365644 374644 365696
rect 374696 365684 374702 365696
rect 379698 365684 379704 365696
rect 374696 365656 379704 365684
rect 374696 365644 374702 365656
rect 379698 365644 379704 365656
rect 379756 365644 379762 365696
rect 539318 365644 539324 365696
rect 539376 365684 539382 365696
rect 542998 365684 543004 365696
rect 539376 365656 543004 365684
rect 539376 365644 539382 365656
rect 542998 365644 543004 365656
rect 543056 365644 543062 365696
rect 211706 365616 211712 365628
rect 190426 365588 211712 365616
rect 211706 365576 211712 365588
rect 211764 365576 211770 365628
rect 222010 365576 222016 365628
rect 222068 365616 222074 365628
rect 232498 365616 232504 365628
rect 222068 365588 232504 365616
rect 222068 365576 222074 365588
rect 232498 365576 232504 365588
rect 232556 365576 232562 365628
rect 249702 365576 249708 365628
rect 249760 365616 249766 365628
rect 260190 365616 260196 365628
rect 249760 365588 260196 365616
rect 249760 365576 249766 365588
rect 260190 365576 260196 365588
rect 260248 365576 260254 365628
rect 261478 365576 261484 365628
rect 261536 365616 261542 365628
rect 567194 365616 567200 365628
rect 261536 365588 567200 365616
rect 261536 365576 261542 365588
rect 567194 365576 567200 365588
rect 567252 365576 567258 365628
rect 53650 365508 53656 365560
rect 53708 365548 53714 365560
rect 69658 365548 69664 365560
rect 53708 365520 69664 365548
rect 53708 365508 53714 365520
rect 69658 365508 69664 365520
rect 69716 365508 69722 365560
rect 81986 365508 81992 365560
rect 82044 365548 82050 365560
rect 94498 365548 94504 365560
rect 82044 365520 94504 365548
rect 82044 365508 82050 365520
rect 94498 365508 94504 365520
rect 94556 365508 94562 365560
rect 109678 365508 109684 365560
rect 109736 365548 109742 365560
rect 120718 365548 120724 365560
rect 109736 365520 120724 365548
rect 109736 365508 109742 365520
rect 120718 365508 120724 365520
rect 120776 365508 120782 365560
rect 137646 365508 137652 365560
rect 137704 365548 137710 365560
rect 148318 365548 148324 365560
rect 137704 365520 148324 365548
rect 137704 365508 137710 365520
rect 148318 365508 148324 365520
rect 148376 365508 148382 365560
rect 193674 365508 193680 365560
rect 193732 365548 193738 365560
rect 204898 365548 204904 365560
rect 193732 365520 204904 365548
rect 193732 365508 193738 365520
rect 204898 365508 204904 365520
rect 204956 365508 204962 365560
rect 238846 365508 238852 365560
rect 238904 365548 238910 365560
rect 268010 365548 268016 365560
rect 238904 365520 268016 365548
rect 238904 365508 238910 365520
rect 268010 365508 268016 365520
rect 268068 365508 268074 365560
rect 277670 365508 277676 365560
rect 277728 365548 277734 365560
rect 289078 365548 289084 365560
rect 277728 365520 289084 365548
rect 277728 365508 277734 365520
rect 289078 365508 289084 365520
rect 289136 365508 289142 365560
rect 306006 365508 306012 365560
rect 306064 365548 306070 365560
rect 316678 365548 316684 365560
rect 306064 365520 316684 365548
rect 306064 365508 306070 365520
rect 316678 365508 316684 365520
rect 316736 365508 316742 365560
rect 323026 365508 323032 365560
rect 323084 365548 323090 365560
rect 352006 365548 352012 365560
rect 323084 365520 352012 365548
rect 323084 365508 323090 365520
rect 352006 365508 352012 365520
rect 352064 365508 352070 365560
rect 361666 365508 361672 365560
rect 361724 365548 361730 365560
rect 373258 365548 373264 365560
rect 361724 365520 373264 365548
rect 361724 365508 361730 365520
rect 373258 365508 373264 365520
rect 373316 365508 373322 365560
rect 379606 365508 379612 365560
rect 379664 365548 379670 365560
rect 408034 365548 408040 365560
rect 379664 365520 408040 365548
rect 379664 365508 379670 365520
rect 408034 365508 408040 365520
rect 408092 365508 408098 365560
rect 417694 365508 417700 365560
rect 417752 365548 417758 365560
rect 428458 365548 428464 365560
rect 417752 365520 428464 365548
rect 417752 365508 417758 365520
rect 428458 365508 428464 365520
rect 428516 365508 428522 365560
rect 434806 365508 434812 365560
rect 434864 365548 434870 365560
rect 463694 365548 463700 365560
rect 434864 365520 463700 365548
rect 434864 365508 434870 365520
rect 463694 365508 463700 365520
rect 463752 365508 463758 365560
rect 473998 365508 474004 365560
rect 474056 365548 474062 365560
rect 485038 365548 485044 365560
rect 474056 365520 485044 365548
rect 474056 365508 474062 365520
rect 485038 365508 485044 365520
rect 485096 365508 485102 365560
rect 501690 365508 501696 365560
rect 501748 365548 501754 365560
rect 512638 365548 512644 365560
rect 501748 365520 512644 365548
rect 501748 365508 501754 365520
rect 512638 365508 512644 365520
rect 512696 365508 512702 365560
rect 518986 365508 518992 365560
rect 519044 365548 519050 365560
rect 547874 365548 547880 365560
rect 519044 365520 547880 365548
rect 519044 365508 519050 365520
rect 547874 365508 547880 365520
rect 547932 365508 547938 365560
rect 333698 365440 333704 365492
rect 333756 365480 333762 365492
rect 344278 365480 344284 365492
rect 333756 365452 344284 365480
rect 333756 365440 333762 365452
rect 344278 365440 344284 365452
rect 344336 365440 344342 365492
rect 390002 365440 390008 365492
rect 390060 365480 390066 365492
rect 400858 365480 400864 365492
rect 390060 365452 400864 365480
rect 390060 365440 390066 365452
rect 400858 365440 400864 365452
rect 400916 365440 400922 365492
rect 445662 365440 445668 365492
rect 445720 365480 445726 365492
rect 456058 365480 456064 365492
rect 445720 365452 456064 365480
rect 445720 365440 445726 365452
rect 456058 365440 456064 365452
rect 456116 365440 456122 365492
rect 529658 365440 529664 365492
rect 529716 365480 529722 365492
rect 540238 365480 540244 365492
rect 529716 365452 540244 365480
rect 529716 365440 529722 365452
rect 540238 365440 540244 365452
rect 540296 365440 540302 365492
rect 36814 365372 36820 365424
rect 36872 365412 36878 365424
rect 557534 365412 557540 365424
rect 36872 365384 557540 365412
rect 36872 365372 36878 365384
rect 557534 365372 557540 365384
rect 557592 365372 557598 365424
rect 16022 362176 16028 362228
rect 16080 362216 16086 362228
rect 547874 362216 547880 362228
rect 16080 362188 547880 362216
rect 16080 362176 16086 362188
rect 547874 362176 547880 362188
rect 547932 362176 547938 362228
rect 25682 361836 25688 361888
rect 25740 361876 25746 361888
rect 261478 361876 261484 361888
rect 25740 361848 261484 361876
rect 25740 361836 25746 361848
rect 261478 361836 261484 361848
rect 261536 361836 261542 361888
rect 148410 361768 148416 361820
rect 148468 361808 148474 361820
rect 165706 361808 165712 361820
rect 148468 361780 165712 361808
rect 148468 361768 148474 361780
rect 165706 361768 165712 361780
rect 165764 361768 165770 361820
rect 175458 361768 175464 361820
rect 175516 361808 175522 361820
rect 193674 361808 193680 361820
rect 175516 361780 193680 361808
rect 175516 361768 175522 361780
rect 193674 361768 193680 361780
rect 193732 361768 193738 361820
rect 203518 361768 203524 361820
rect 203576 361808 203582 361820
rect 221366 361808 221372 361820
rect 203576 361780 221372 361808
rect 203576 361768 203582 361780
rect 221366 361768 221372 361780
rect 221424 361768 221430 361820
rect 296346 361768 296352 361820
rect 296404 361808 296410 361820
rect 316770 361808 316776 361820
rect 296404 361780 316776 361808
rect 296404 361768 296410 361780
rect 316770 361768 316776 361780
rect 316828 361768 316834 361820
rect 408034 361768 408040 361820
rect 408092 361808 408098 361820
rect 428642 361808 428648 361820
rect 408092 361780 428648 361808
rect 408092 361768 408098 361780
rect 428642 361768 428648 361780
rect 428700 361768 428706 361820
rect 492030 361768 492036 361820
rect 492088 361808 492094 361820
rect 512730 361808 512736 361820
rect 492088 361780 512736 361808
rect 492088 361768 492094 361780
rect 512730 361768 512736 361780
rect 512788 361768 512794 361820
rect 36998 361700 37004 361752
rect 37056 361740 37062 361752
rect 53650 361740 53656 361752
rect 37056 361712 53656 361740
rect 37056 361700 37062 361712
rect 53650 361700 53656 361712
rect 53708 361700 53714 361752
rect 64322 361700 64328 361752
rect 64380 361740 64386 361752
rect 81434 361740 81440 361752
rect 64380 361712 81440 361740
rect 64380 361700 64386 361712
rect 81434 361700 81440 361712
rect 81492 361700 81498 361752
rect 91462 361700 91468 361752
rect 91520 361740 91526 361752
rect 109678 361740 109684 361752
rect 91520 361712 109684 361740
rect 91520 361700 91526 361712
rect 109678 361700 109684 361712
rect 109736 361700 109742 361752
rect 119430 361700 119436 361752
rect 119488 361740 119494 361752
rect 137646 361740 137652 361752
rect 119488 361712 137652 361740
rect 119488 361700 119494 361712
rect 137646 361700 137652 361712
rect 137704 361700 137710 361752
rect 156322 361700 156328 361752
rect 156380 361740 156386 361752
rect 178678 361740 178684 361752
rect 156380 361712 178684 361740
rect 156380 361700 156386 361712
rect 178678 361700 178684 361712
rect 178736 361700 178742 361752
rect 232590 361700 232596 361752
rect 232648 361740 232654 361752
rect 249702 361740 249708 361752
rect 232648 361712 249708 361740
rect 232648 361700 232654 361712
rect 249702 361700 249708 361712
rect 249760 361700 249766 361752
rect 260098 361700 260104 361752
rect 260156 361740 260162 361752
rect 277670 361740 277676 361752
rect 260156 361712 277676 361740
rect 260156 361700 260162 361712
rect 277670 361700 277676 361712
rect 277728 361700 277734 361752
rect 287514 361700 287520 361752
rect 287572 361740 287578 361752
rect 305362 361740 305368 361752
rect 287572 361712 305368 361740
rect 287572 361700 287578 361712
rect 305362 361700 305368 361712
rect 305420 361700 305426 361752
rect 345658 361700 345664 361752
rect 345716 361740 345722 361752
rect 361666 361740 361672 361752
rect 345716 361712 361672 361740
rect 345716 361700 345722 361712
rect 361666 361700 361672 361712
rect 361724 361700 361730 361752
rect 371510 361700 371516 361752
rect 371568 361740 371574 361752
rect 389358 361740 389364 361752
rect 371568 361712 389364 361740
rect 371568 361700 371574 361712
rect 389358 361700 389364 361712
rect 389416 361700 389422 361752
rect 399478 361700 399484 361752
rect 399536 361740 399542 361752
rect 417694 361740 417700 361752
rect 399536 361712 417700 361740
rect 399536 361700 399542 361712
rect 417694 361700 417700 361712
rect 417752 361700 417758 361752
rect 456058 361700 456064 361752
rect 456116 361740 456122 361752
rect 473354 361740 473360 361752
rect 456116 361712 473360 361740
rect 456116 361700 456122 361712
rect 473354 361700 473360 361712
rect 473412 361700 473418 361752
rect 483474 361700 483480 361752
rect 483532 361740 483538 361752
rect 501690 361740 501696 361752
rect 483532 361712 501696 361740
rect 483532 361700 483538 361712
rect 501690 361700 501696 361712
rect 501748 361700 501754 361752
rect 36814 361632 36820 361684
rect 36872 361672 36878 361684
rect 63310 361672 63316 361684
rect 36872 361644 63316 361672
rect 36872 361632 36878 361644
rect 63310 361632 63316 361644
rect 63368 361632 63374 361684
rect 66898 361632 66904 361684
rect 66956 361672 66962 361684
rect 91094 361672 91100 361684
rect 66956 361644 91100 361672
rect 66956 361632 66962 361644
rect 91094 361632 91100 361644
rect 91152 361632 91158 361684
rect 94498 361632 94504 361684
rect 94556 361672 94562 361684
rect 119338 361672 119344 361684
rect 94556 361644 119344 361672
rect 94556 361632 94562 361644
rect 119338 361632 119344 361644
rect 119396 361632 119402 361684
rect 120718 361632 120724 361684
rect 120776 361672 120782 361684
rect 147306 361672 147312 361684
rect 120776 361644 147312 361672
rect 120776 361632 120782 361644
rect 147306 361632 147312 361644
rect 147364 361632 147370 361684
rect 148318 361632 148324 361684
rect 148376 361672 148382 361684
rect 175366 361672 175372 361684
rect 148376 361644 175372 361672
rect 148376 361632 148382 361644
rect 175366 361632 175372 361644
rect 175424 361632 175430 361684
rect 177298 361632 177304 361684
rect 177356 361672 177362 361684
rect 203334 361672 203340 361684
rect 177356 361644 203340 361672
rect 177356 361632 177362 361644
rect 203334 361632 203340 361644
rect 203392 361632 203398 361684
rect 204898 361632 204904 361684
rect 204956 361672 204962 361684
rect 231026 361672 231032 361684
rect 204956 361644 231032 361672
rect 204956 361632 204962 361644
rect 231026 361632 231032 361644
rect 231084 361632 231090 361684
rect 232498 361632 232504 361684
rect 232556 361672 232562 361684
rect 259362 361672 259368 361684
rect 232556 361644 259368 361672
rect 232556 361632 232562 361644
rect 259362 361632 259368 361644
rect 259420 361632 259426 361684
rect 268010 361632 268016 361684
rect 268068 361672 268074 361684
rect 287698 361672 287704 361684
rect 268068 361644 287704 361672
rect 268068 361632 268074 361644
rect 287698 361632 287704 361644
rect 287756 361632 287762 361684
rect 315482 361632 315488 361684
rect 315540 361672 315546 361684
rect 333698 361672 333704 361684
rect 315540 361644 333704 361672
rect 315540 361632 315546 361644
rect 333698 361632 333704 361644
rect 333756 361632 333762 361684
rect 352006 361632 352012 361684
rect 352064 361672 352070 361684
rect 374638 361672 374644 361684
rect 352064 361644 374644 361672
rect 352064 361632 352070 361644
rect 374638 361632 374644 361644
rect 374696 361632 374702 361684
rect 428550 361632 428556 361684
rect 428608 361672 428614 361684
rect 445662 361672 445668 361684
rect 428608 361644 445668 361672
rect 428608 361632 428614 361644
rect 445662 361632 445668 361644
rect 445720 361632 445726 361684
rect 464338 361632 464344 361684
rect 464396 361672 464402 361684
rect 483658 361672 483664 361684
rect 464396 361644 483664 361672
rect 464396 361632 464402 361644
rect 483658 361632 483664 361644
rect 483716 361632 483722 361684
rect 511442 361632 511448 361684
rect 511500 361672 511506 361684
rect 529658 361672 529664 361684
rect 511500 361644 529664 361672
rect 511500 361632 511506 361644
rect 529658 361632 529664 361644
rect 529716 361632 529722 361684
rect 542998 361632 543004 361684
rect 543056 361672 543062 361684
rect 557534 361672 557540 361684
rect 543056 361644 557540 361672
rect 543056 361632 543062 361644
rect 557534 361632 557540 361644
rect 557592 361632 557598 361684
rect 212350 361564 212356 361616
rect 212408 361604 212414 361616
rect 232682 361604 232688 361616
rect 212408 361576 232688 361604
rect 212408 361564 212414 361576
rect 232682 361564 232688 361576
rect 232740 361564 232746 361616
rect 260190 361564 260196 361616
rect 260248 361604 260254 361616
rect 287330 361604 287336 361616
rect 260248 361576 287336 361604
rect 260248 361564 260254 361576
rect 287330 361564 287336 361576
rect 287388 361564 287394 361616
rect 289078 361564 289084 361616
rect 289136 361604 289142 361616
rect 315022 361604 315028 361616
rect 289136 361576 315028 361604
rect 289136 361564 289142 361576
rect 315022 361564 315028 361576
rect 315080 361564 315086 361616
rect 316678 361564 316684 361616
rect 316736 361604 316742 361616
rect 343358 361604 343364 361616
rect 316736 361576 343364 361604
rect 316736 361564 316742 361576
rect 343358 361564 343364 361576
rect 343416 361564 343422 361616
rect 344278 361564 344284 361616
rect 344336 361604 344342 361616
rect 371326 361604 371332 361616
rect 344336 361576 371332 361604
rect 344336 361564 344342 361576
rect 371326 361564 371332 361576
rect 371384 361564 371390 361616
rect 373258 361564 373264 361616
rect 373316 361604 373322 361616
rect 399018 361604 399024 361616
rect 373316 361576 399024 361604
rect 373316 361564 373322 361576
rect 399018 361564 399024 361576
rect 399076 361564 399082 361616
rect 400858 361564 400864 361616
rect 400916 361604 400922 361616
rect 427354 361604 427360 361616
rect 400916 361576 427360 361604
rect 400916 361564 400922 361576
rect 427354 361564 427360 361576
rect 427412 361564 427418 361616
rect 428458 361564 428464 361616
rect 428516 361604 428522 361616
rect 455322 361604 455328 361616
rect 428516 361576 455328 361604
rect 428516 361564 428522 361576
rect 455322 361564 455328 361576
rect 455380 361564 455386 361616
rect 456150 361564 456156 361616
rect 456208 361604 456214 361616
rect 483014 361604 483020 361616
rect 456208 361576 483020 361604
rect 456208 361564 456214 361576
rect 483014 361564 483020 361576
rect 483072 361564 483078 361616
rect 485038 361564 485044 361616
rect 485096 361604 485102 361616
rect 511350 361604 511356 361616
rect 485096 361576 511356 361604
rect 485096 361564 485102 361576
rect 511350 361564 511356 361576
rect 511408 361564 511414 361616
rect 512638 361564 512644 361616
rect 512696 361604 512702 361616
rect 539318 361604 539324 361616
rect 512696 361576 539324 361604
rect 512696 361564 512702 361576
rect 539318 361564 539324 361576
rect 539376 361564 539382 361616
rect 540238 361564 540244 361616
rect 540296 361604 540302 361616
rect 567194 361604 567200 361616
rect 540296 361576 567200 361604
rect 540296 361564 540302 361576
rect 567194 361564 567200 361576
rect 567252 361564 567258 361616
rect 37918 359456 37924 359508
rect 37976 359496 37982 359508
rect 545758 359496 545764 359508
rect 37976 359468 545764 359496
rect 37976 359456 37982 359468
rect 545758 359456 545764 359468
rect 545816 359456 545822 359508
rect 35618 358776 35624 358828
rect 35676 358816 35682 358828
rect 36906 358816 36912 358828
rect 35676 358788 36912 358816
rect 35676 358776 35682 358788
rect 36906 358776 36912 358788
rect 36964 358776 36970 358828
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 14458 357456 14464 357468
rect 3384 357428 14464 357456
rect 3384 357416 3390 357428
rect 14458 357416 14464 357428
rect 14516 357416 14522 357468
rect 63586 342524 63592 342576
rect 63644 342564 63650 342576
rect 64322 342564 64328 342576
rect 63644 342536 64328 342564
rect 63644 342524 63650 342536
rect 64322 342524 64328 342536
rect 64380 342524 64386 342576
rect 147674 342524 147680 342576
rect 147732 342564 147738 342576
rect 148410 342564 148416 342576
rect 147732 342536 148416 342564
rect 147732 342524 147738 342536
rect 148410 342524 148416 342536
rect 148468 342524 148474 342576
rect 316770 341912 316776 341964
rect 316828 341952 316834 341964
rect 323670 341952 323676 341964
rect 316828 341924 323676 341952
rect 316828 341912 316834 341924
rect 323670 341912 323676 341924
rect 323728 341912 323734 341964
rect 512730 341912 512736 341964
rect 512788 341952 512794 341964
rect 519630 341952 519636 341964
rect 512788 341924 519636 341952
rect 512788 341912 512794 341924
rect 519630 341912 519636 341924
rect 519688 341912 519694 341964
rect 287698 341504 287704 341556
rect 287756 341544 287762 341556
rect 295702 341544 295708 341556
rect 287756 341516 295708 341544
rect 287756 341504 287762 341516
rect 295702 341504 295708 341516
rect 295760 341504 295766 341556
rect 428642 341504 428648 341556
rect 428700 341544 428706 341556
rect 435726 341544 435732 341556
rect 428700 341516 435732 341544
rect 428700 341504 428706 341516
rect 435726 341504 435732 341516
rect 435784 341504 435790 341556
rect 232682 341368 232688 341420
rect 232740 341408 232746 341420
rect 239766 341408 239772 341420
rect 232740 341380 239772 341408
rect 232740 341368 232746 341380
rect 239766 341368 239772 341380
rect 239824 341368 239830 341420
rect 483658 341368 483664 341420
rect 483716 341408 483722 341420
rect 491662 341408 491668 341420
rect 483716 341380 491668 341408
rect 483716 341368 483722 341380
rect 491662 341368 491668 341380
rect 491720 341368 491726 341420
rect 13722 340824 13728 340876
rect 13780 340864 13786 340876
rect 66254 340864 66260 340876
rect 13780 340836 66260 340864
rect 13780 340824 13786 340836
rect 66254 340824 66260 340836
rect 66312 340824 66318 340876
rect 70302 340824 70308 340876
rect 70360 340864 70366 340876
rect 121454 340864 121460 340876
rect 70360 340836 121460 340864
rect 70360 340824 70366 340836
rect 121454 340824 121460 340836
rect 121512 340824 121518 340876
rect 126882 340824 126888 340876
rect 126940 340864 126946 340876
rect 178034 340864 178040 340876
rect 126940 340836 178040 340864
rect 126940 340824 126946 340836
rect 178034 340824 178040 340836
rect 178092 340824 178098 340876
rect 209682 340824 209688 340876
rect 209740 340864 209746 340876
rect 262214 340864 262220 340876
rect 209740 340836 262220 340864
rect 209740 340824 209746 340836
rect 262214 340824 262220 340836
rect 262272 340824 262278 340876
rect 266262 340824 266268 340876
rect 266320 340864 266326 340876
rect 317414 340864 317420 340876
rect 266320 340836 317420 340864
rect 266320 340824 266326 340836
rect 317414 340824 317420 340836
rect 317472 340824 317478 340876
rect 322842 340824 322848 340876
rect 322900 340864 322906 340876
rect 373994 340864 374000 340876
rect 322900 340836 374000 340864
rect 322900 340824 322906 340836
rect 373994 340824 374000 340836
rect 374052 340824 374058 340876
rect 405642 340824 405648 340876
rect 405700 340864 405706 340876
rect 458174 340864 458180 340876
rect 405700 340836 458180 340864
rect 405700 340824 405706 340836
rect 458174 340824 458180 340836
rect 458232 340824 458238 340876
rect 489822 340824 489828 340876
rect 489880 340864 489886 340876
rect 542354 340864 542360 340876
rect 489880 340836 542360 340864
rect 489880 340824 489886 340836
rect 542354 340824 542360 340836
rect 542412 340824 542418 340876
rect 35618 340756 35624 340808
rect 35676 340796 35682 340808
rect 36998 340796 37004 340808
rect 35676 340768 37004 340796
rect 35676 340756 35682 340768
rect 36998 340756 37004 340768
rect 37056 340756 37062 340808
rect 42702 340756 42708 340808
rect 42760 340796 42766 340808
rect 93854 340796 93860 340808
rect 42760 340768 93860 340796
rect 42760 340756 42766 340768
rect 93854 340756 93860 340768
rect 93912 340756 93918 340808
rect 97902 340756 97908 340808
rect 97960 340796 97966 340808
rect 149054 340796 149060 340808
rect 97960 340768 149060 340796
rect 97960 340756 97966 340768
rect 149054 340756 149060 340768
rect 149112 340756 149118 340808
rect 154482 340756 154488 340808
rect 154540 340796 154546 340808
rect 205634 340796 205640 340808
rect 154540 340768 205640 340796
rect 154540 340756 154546 340768
rect 205634 340756 205640 340768
rect 205692 340756 205698 340808
rect 231670 340756 231676 340808
rect 231728 340796 231734 340808
rect 232590 340796 232596 340808
rect 231728 340768 232596 340796
rect 231728 340756 231734 340768
rect 232590 340756 232596 340768
rect 232648 340756 232654 340808
rect 238662 340756 238668 340808
rect 238720 340796 238726 340808
rect 289814 340796 289820 340808
rect 238720 340768 289820 340796
rect 238720 340756 238726 340768
rect 289814 340756 289820 340768
rect 289872 340756 289878 340808
rect 293862 340756 293868 340808
rect 293920 340796 293926 340808
rect 345014 340796 345020 340808
rect 293920 340768 345020 340796
rect 293920 340756 293926 340768
rect 345014 340756 345020 340768
rect 345072 340756 345078 340808
rect 350442 340756 350448 340808
rect 350500 340796 350506 340808
rect 401594 340796 401600 340808
rect 350500 340768 401600 340796
rect 350500 340756 350506 340768
rect 401594 340756 401600 340768
rect 401652 340756 401658 340808
rect 427722 340756 427728 340808
rect 427780 340796 427786 340808
rect 428550 340796 428556 340808
rect 427780 340768 428556 340796
rect 427780 340756 427786 340768
rect 428550 340756 428556 340768
rect 428608 340756 428614 340808
rect 434622 340756 434628 340808
rect 434680 340796 434686 340808
rect 485774 340796 485780 340808
rect 434680 340768 485780 340796
rect 434680 340756 434686 340768
rect 485774 340756 485780 340768
rect 485832 340756 485838 340808
rect 518802 340756 518808 340808
rect 518860 340796 518866 340808
rect 569954 340796 569960 340808
rect 518860 340768 569960 340796
rect 518860 340756 518866 340768
rect 569954 340756 569960 340768
rect 570012 340756 570018 340808
rect 182082 340688 182088 340740
rect 182140 340728 182146 340740
rect 233234 340728 233240 340740
rect 182140 340700 233240 340728
rect 182140 340688 182146 340700
rect 233234 340688 233240 340700
rect 233292 340688 233298 340740
rect 343634 340688 343640 340740
rect 343692 340728 343698 340740
rect 345658 340728 345664 340740
rect 343692 340700 345664 340728
rect 343692 340688 343698 340700
rect 345658 340688 345664 340700
rect 345716 340688 345722 340740
rect 378042 340688 378048 340740
rect 378100 340728 378106 340740
rect 429194 340728 429200 340740
rect 378100 340700 429200 340728
rect 378100 340688 378106 340700
rect 429194 340688 429200 340700
rect 429252 340688 429258 340740
rect 462222 340688 462228 340740
rect 462280 340728 462286 340740
rect 513374 340728 513380 340740
rect 462280 340700 513380 340728
rect 462280 340688 462286 340700
rect 513374 340688 513380 340700
rect 513432 340688 513438 340740
rect 539502 340688 539508 340740
rect 539560 340728 539566 340740
rect 542998 340728 543004 340740
rect 539560 340700 543004 340728
rect 539560 340688 539566 340700
rect 542998 340688 543004 340700
rect 543056 340688 543062 340740
rect 178678 338036 178684 338088
rect 178736 338076 178742 338088
rect 184014 338076 184020 338088
rect 178736 338048 184020 338076
rect 178736 338036 178742 338048
rect 184014 338036 184020 338048
rect 184072 338036 184078 338088
rect 374638 338036 374644 338088
rect 374696 338076 374702 338088
rect 379698 338076 379704 338088
rect 374696 338048 379704 338076
rect 374696 338036 374702 338048
rect 379698 338036 379704 338048
rect 379756 338036 379762 338088
rect 15194 337968 15200 338020
rect 15252 338008 15258 338020
rect 43990 338008 43996 338020
rect 15252 337980 43996 338008
rect 15252 337968 15258 337980
rect 43990 337968 43996 337980
rect 44048 337968 44054 338020
rect 71038 337968 71044 338020
rect 71096 338008 71102 338020
rect 567194 338008 567200 338020
rect 71096 337980 567200 338008
rect 71096 337968 71102 337980
rect 567194 337968 567200 337980
rect 567252 337968 567258 338020
rect 25682 337900 25688 337952
rect 25740 337940 25746 337952
rect 36814 337940 36820 337952
rect 25740 337912 36820 337940
rect 25740 337900 25746 337912
rect 36814 337900 36820 337912
rect 36872 337900 36878 337952
rect 53650 337900 53656 337952
rect 53708 337940 53714 337952
rect 66898 337940 66904 337952
rect 53708 337912 66904 337940
rect 53708 337900 53714 337912
rect 66898 337900 66904 337912
rect 66956 337900 66962 337952
rect 71866 337900 71872 337952
rect 71924 337940 71930 337952
rect 100018 337940 100024 337952
rect 71924 337912 100024 337940
rect 71924 337900 71930 337912
rect 100018 337900 100024 337912
rect 100076 337900 100082 337952
rect 127986 337940 127992 337952
rect 103486 337912 127992 337940
rect 42886 337832 42892 337884
rect 42944 337872 42950 337884
rect 72050 337872 72056 337884
rect 42944 337844 72056 337872
rect 42944 337832 42950 337844
rect 72050 337832 72056 337844
rect 72108 337832 72114 337884
rect 81986 337832 81992 337884
rect 82044 337872 82050 337884
rect 94498 337872 94504 337884
rect 82044 337844 94504 337872
rect 82044 337832 82050 337844
rect 94498 337832 94504 337844
rect 94556 337832 94562 337884
rect 99466 337832 99472 337884
rect 99524 337872 99530 337884
rect 103486 337872 103514 337912
rect 127986 337900 127992 337912
rect 128044 337900 128050 337952
rect 156046 337940 156052 337952
rect 132466 337912 156052 337940
rect 99524 337844 103514 337872
rect 99524 337832 99530 337844
rect 109678 337832 109684 337884
rect 109736 337872 109742 337884
rect 120718 337872 120724 337884
rect 109736 337844 120724 337872
rect 109736 337832 109742 337844
rect 120718 337832 120724 337844
rect 120776 337832 120782 337884
rect 127066 337832 127072 337884
rect 127124 337872 127130 337884
rect 132466 337872 132494 337912
rect 156046 337900 156052 337912
rect 156104 337900 156110 337952
rect 165982 337900 165988 337952
rect 166040 337940 166046 337952
rect 177298 337940 177304 337952
rect 166040 337912 177304 337940
rect 166040 337900 166046 337912
rect 177298 337900 177304 337912
rect 177356 337900 177362 337952
rect 183646 337900 183652 337952
rect 183704 337940 183710 337952
rect 211706 337940 211712 337952
rect 183704 337912 211712 337940
rect 183704 337900 183710 337912
rect 211706 337900 211712 337912
rect 211764 337900 211770 337952
rect 222010 337900 222016 337952
rect 222068 337940 222074 337952
rect 232498 337940 232504 337952
rect 222068 337912 232504 337940
rect 222068 337900 222074 337912
rect 232498 337900 232504 337912
rect 232556 337900 232562 337952
rect 238846 337900 238852 337952
rect 238904 337940 238910 337952
rect 268010 337940 268016 337952
rect 238904 337912 268016 337940
rect 238904 337900 238910 337912
rect 268010 337900 268016 337912
rect 268068 337900 268074 337952
rect 277670 337900 277676 337952
rect 277728 337940 277734 337952
rect 289078 337940 289084 337952
rect 277728 337912 289084 337940
rect 277728 337900 277734 337912
rect 289078 337900 289084 337912
rect 289136 337900 289142 337952
rect 306006 337900 306012 337952
rect 306064 337940 306070 337952
rect 316678 337940 316684 337952
rect 306064 337912 316684 337940
rect 306064 337900 306070 337912
rect 316678 337900 316684 337912
rect 316736 337900 316742 337952
rect 323026 337900 323032 337952
rect 323084 337940 323090 337952
rect 352006 337940 352012 337952
rect 323084 337912 352012 337940
rect 323084 337900 323090 337912
rect 352006 337900 352012 337912
rect 352064 337900 352070 337952
rect 361666 337900 361672 337952
rect 361724 337940 361730 337952
rect 373258 337940 373264 337952
rect 361724 337912 373264 337940
rect 361724 337900 361730 337912
rect 373258 337900 373264 337912
rect 373316 337900 373322 337952
rect 379606 337900 379612 337952
rect 379664 337940 379670 337952
rect 408034 337940 408040 337952
rect 379664 337912 408040 337940
rect 379664 337900 379670 337912
rect 408034 337900 408040 337912
rect 408092 337900 408098 337952
rect 417694 337900 417700 337952
rect 417752 337940 417758 337952
rect 428458 337940 428464 337952
rect 417752 337912 428464 337940
rect 417752 337900 417758 337912
rect 428458 337900 428464 337912
rect 428516 337900 428522 337952
rect 434806 337900 434812 337952
rect 434864 337940 434870 337952
rect 463694 337940 463700 337952
rect 434864 337912 463700 337940
rect 434864 337900 434870 337912
rect 463694 337900 463700 337912
rect 463752 337900 463758 337952
rect 473998 337900 474004 337952
rect 474056 337940 474062 337952
rect 485038 337940 485044 337952
rect 474056 337912 485044 337940
rect 474056 337900 474062 337912
rect 485038 337900 485044 337912
rect 485096 337900 485102 337952
rect 501690 337900 501696 337952
rect 501748 337940 501754 337952
rect 512638 337940 512644 337952
rect 501748 337912 512644 337940
rect 501748 337900 501754 337912
rect 512638 337900 512644 337912
rect 512696 337900 512702 337952
rect 518986 337900 518992 337952
rect 519044 337940 519050 337952
rect 547874 337940 547880 337952
rect 519044 337912 547880 337940
rect 519044 337900 519050 337912
rect 547874 337900 547880 337912
rect 547932 337900 547938 337952
rect 127124 337844 132494 337872
rect 127124 337832 127130 337844
rect 137646 337832 137652 337884
rect 137704 337872 137710 337884
rect 148318 337872 148324 337884
rect 137704 337844 148324 337872
rect 137704 337832 137710 337844
rect 148318 337832 148324 337844
rect 148376 337832 148382 337884
rect 193674 337832 193680 337884
rect 193732 337872 193738 337884
rect 204898 337872 204904 337884
rect 193732 337844 204904 337872
rect 193732 337832 193738 337844
rect 204898 337832 204904 337844
rect 204956 337832 204962 337884
rect 249702 337832 249708 337884
rect 249760 337872 249766 337884
rect 260190 337872 260196 337884
rect 249760 337844 260196 337872
rect 249760 337832 249766 337844
rect 260190 337832 260196 337844
rect 260248 337832 260254 337884
rect 333698 337832 333704 337884
rect 333756 337872 333762 337884
rect 344278 337872 344284 337884
rect 333756 337844 344284 337872
rect 333756 337832 333762 337844
rect 344278 337832 344284 337844
rect 344336 337832 344342 337884
rect 390002 337832 390008 337884
rect 390060 337872 390066 337884
rect 400858 337872 400864 337884
rect 390060 337844 400864 337872
rect 390060 337832 390066 337844
rect 400858 337832 400864 337844
rect 400916 337832 400922 337884
rect 445662 337832 445668 337884
rect 445720 337872 445726 337884
rect 456150 337872 456156 337884
rect 445720 337844 456156 337872
rect 445720 337832 445726 337844
rect 456150 337832 456156 337844
rect 456208 337832 456214 337884
rect 529658 337832 529664 337884
rect 529716 337872 529722 337884
rect 540238 337872 540244 337884
rect 529716 337844 540244 337872
rect 529716 337832 529722 337844
rect 540238 337832 540244 337844
rect 540296 337832 540302 337884
rect 36722 337764 36728 337816
rect 36780 337804 36786 337816
rect 557534 337804 557540 337816
rect 36780 337776 557540 337804
rect 36780 337764 36786 337776
rect 557534 337764 557540 337776
rect 557592 337764 557598 337816
rect 16022 335996 16028 336048
rect 16080 336036 16086 336048
rect 547874 336036 547880 336048
rect 16080 336008 547880 336036
rect 16080 335996 16086 336008
rect 547874 335996 547880 336008
rect 547932 335996 547938 336048
rect 25682 335520 25688 335572
rect 25740 335560 25746 335572
rect 71038 335560 71044 335572
rect 25740 335532 71044 335560
rect 25740 335520 25746 335532
rect 71038 335520 71044 335532
rect 71096 335520 71102 335572
rect 212258 335520 212264 335572
rect 212316 335560 212322 335572
rect 232682 335560 232688 335572
rect 212316 335532 232688 335560
rect 212316 335520 212322 335532
rect 232682 335520 232688 335532
rect 232740 335520 232746 335572
rect 296346 335520 296352 335572
rect 296404 335560 296410 335572
rect 316770 335560 316776 335572
rect 296404 335532 316776 335560
rect 296404 335520 296410 335532
rect 316770 335520 316776 335532
rect 316828 335520 316834 335572
rect 408034 335520 408040 335572
rect 408092 335560 408098 335572
rect 428642 335560 428648 335572
rect 408092 335532 428648 335560
rect 408092 335520 408098 335532
rect 428642 335520 428648 335532
rect 428700 335520 428706 335572
rect 492030 335520 492036 335572
rect 492088 335560 492094 335572
rect 512730 335560 512736 335572
rect 492088 335532 512736 335560
rect 492088 335520 492094 335532
rect 512730 335520 512736 335532
rect 512788 335520 512794 335572
rect 36998 335452 37004 335504
rect 37056 335492 37062 335504
rect 53650 335492 53656 335504
rect 37056 335464 53656 335492
rect 37056 335452 37062 335464
rect 53650 335452 53656 335464
rect 53708 335452 53714 335504
rect 148318 335452 148324 335504
rect 148376 335492 148382 335504
rect 165614 335492 165620 335504
rect 148376 335464 165620 335492
rect 148376 335452 148382 335464
rect 165614 335452 165620 335464
rect 165672 335452 165678 335504
rect 175458 335452 175464 335504
rect 175516 335492 175522 335504
rect 193674 335492 193680 335504
rect 175516 335464 193680 335492
rect 175516 335452 175522 335464
rect 193674 335452 193680 335464
rect 193732 335452 193738 335504
rect 203518 335452 203524 335504
rect 203576 335492 203582 335504
rect 221366 335492 221372 335504
rect 203576 335464 221372 335492
rect 203576 335452 203582 335464
rect 221366 335452 221372 335464
rect 221424 335452 221430 335504
rect 260190 335452 260196 335504
rect 260248 335492 260254 335504
rect 277670 335492 277676 335504
rect 260248 335464 277676 335492
rect 260248 335452 260254 335464
rect 277670 335452 277676 335464
rect 277728 335452 277734 335504
rect 287514 335452 287520 335504
rect 287572 335492 287578 335504
rect 305362 335492 305368 335504
rect 287572 335464 305368 335492
rect 287572 335452 287578 335464
rect 305362 335452 305368 335464
rect 305420 335452 305426 335504
rect 345658 335452 345664 335504
rect 345716 335492 345722 335504
rect 361666 335492 361672 335504
rect 345716 335464 361672 335492
rect 345716 335452 345722 335464
rect 361666 335452 361672 335464
rect 361724 335452 361730 335504
rect 371510 335452 371516 335504
rect 371568 335492 371574 335504
rect 389358 335492 389364 335504
rect 371568 335464 389364 335492
rect 371568 335452 371574 335464
rect 389358 335452 389364 335464
rect 389416 335452 389422 335504
rect 399478 335452 399484 335504
rect 399536 335492 399542 335504
rect 417694 335492 417700 335504
rect 399536 335464 417700 335492
rect 399536 335452 399542 335464
rect 417694 335452 417700 335464
rect 417752 335452 417758 335504
rect 456150 335452 456156 335504
rect 456208 335492 456214 335504
rect 473538 335492 473544 335504
rect 456208 335464 473544 335492
rect 456208 335452 456214 335464
rect 473538 335452 473544 335464
rect 473596 335452 473602 335504
rect 483474 335452 483480 335504
rect 483532 335492 483538 335504
rect 501690 335492 501696 335504
rect 483532 335464 501696 335492
rect 483532 335452 483538 335464
rect 501690 335452 501696 335464
rect 501748 335452 501754 335504
rect 36722 335384 36728 335436
rect 36780 335424 36786 335436
rect 63310 335424 63316 335436
rect 36780 335396 63316 335424
rect 36780 335384 36786 335396
rect 63310 335384 63316 335396
rect 63368 335384 63374 335436
rect 64322 335384 64328 335436
rect 64380 335424 64386 335436
rect 81434 335424 81440 335436
rect 64380 335396 81440 335424
rect 64380 335384 64386 335396
rect 81434 335384 81440 335396
rect 81492 335384 81498 335436
rect 91462 335384 91468 335436
rect 91520 335424 91526 335436
rect 109678 335424 109684 335436
rect 91520 335396 109684 335424
rect 91520 335384 91526 335396
rect 109678 335384 109684 335396
rect 109736 335384 109742 335436
rect 119430 335384 119436 335436
rect 119488 335424 119494 335436
rect 137646 335424 137652 335436
rect 119488 335396 137652 335424
rect 119488 335384 119494 335396
rect 137646 335384 137652 335396
rect 137704 335384 137710 335436
rect 156322 335384 156328 335436
rect 156380 335424 156386 335436
rect 178678 335424 178684 335436
rect 156380 335396 178684 335424
rect 156380 335384 156386 335396
rect 178678 335384 178684 335396
rect 178736 335384 178742 335436
rect 232498 335384 232504 335436
rect 232556 335424 232562 335436
rect 249702 335424 249708 335436
rect 232556 335396 249708 335424
rect 232556 335384 232562 335396
rect 249702 335384 249708 335396
rect 249760 335384 249766 335436
rect 268010 335384 268016 335436
rect 268068 335424 268074 335436
rect 287698 335424 287704 335436
rect 268068 335396 287704 335424
rect 268068 335384 268074 335396
rect 287698 335384 287704 335396
rect 287756 335384 287762 335436
rect 315482 335384 315488 335436
rect 315540 335424 315546 335436
rect 333698 335424 333704 335436
rect 315540 335396 333704 335424
rect 315540 335384 315546 335396
rect 333698 335384 333704 335396
rect 333756 335384 333762 335436
rect 352006 335384 352012 335436
rect 352064 335424 352070 335436
rect 374638 335424 374644 335436
rect 352064 335396 374644 335424
rect 352064 335384 352070 335396
rect 374638 335384 374644 335396
rect 374696 335384 374702 335436
rect 428550 335384 428556 335436
rect 428608 335424 428614 335436
rect 445662 335424 445668 335436
rect 428608 335396 445668 335424
rect 428608 335384 428614 335396
rect 445662 335384 445668 335396
rect 445720 335384 445726 335436
rect 464338 335384 464344 335436
rect 464396 335424 464402 335436
rect 483658 335424 483664 335436
rect 464396 335396 483664 335424
rect 464396 335384 464402 335396
rect 483658 335384 483664 335396
rect 483716 335384 483722 335436
rect 511442 335384 511448 335436
rect 511500 335424 511506 335436
rect 529658 335424 529664 335436
rect 511500 335396 529664 335424
rect 511500 335384 511506 335396
rect 529658 335384 529664 335396
rect 529716 335384 529722 335436
rect 542998 335384 543004 335436
rect 543056 335424 543062 335436
rect 557534 335424 557540 335436
rect 543056 335396 557540 335424
rect 543056 335384 543062 335396
rect 557534 335384 557540 335396
rect 557592 335384 557598 335436
rect 69658 335316 69664 335368
rect 69716 335356 69722 335368
rect 91094 335356 91100 335368
rect 69716 335328 91100 335356
rect 69716 335316 69722 335328
rect 91094 335316 91100 335328
rect 91152 335316 91158 335368
rect 94498 335316 94504 335368
rect 94556 335356 94562 335368
rect 119338 335356 119344 335368
rect 94556 335328 119344 335356
rect 94556 335316 94562 335328
rect 119338 335316 119344 335328
rect 119396 335316 119402 335368
rect 120718 335316 120724 335368
rect 120776 335356 120782 335368
rect 147306 335356 147312 335368
rect 120776 335328 147312 335356
rect 120776 335316 120782 335328
rect 147306 335316 147312 335328
rect 147364 335316 147370 335368
rect 148410 335316 148416 335368
rect 148468 335356 148474 335368
rect 175274 335356 175280 335368
rect 148468 335328 175280 335356
rect 148468 335316 148474 335328
rect 175274 335316 175280 335328
rect 175332 335316 175338 335368
rect 177298 335316 177304 335368
rect 177356 335356 177362 335368
rect 203334 335356 203340 335368
rect 177356 335328 203340 335356
rect 177356 335316 177362 335328
rect 203334 335316 203340 335328
rect 203392 335316 203398 335368
rect 204898 335316 204904 335368
rect 204956 335356 204962 335368
rect 231026 335356 231032 335368
rect 204956 335328 231032 335356
rect 204956 335316 204962 335328
rect 231026 335316 231032 335328
rect 231084 335316 231090 335368
rect 232590 335316 232596 335368
rect 232648 335356 232654 335368
rect 259362 335356 259368 335368
rect 232648 335328 259368 335356
rect 232648 335316 232654 335328
rect 259362 335316 259368 335328
rect 259420 335316 259426 335368
rect 260098 335316 260104 335368
rect 260156 335356 260162 335368
rect 287330 335356 287336 335368
rect 260156 335328 287336 335356
rect 260156 335316 260162 335328
rect 287330 335316 287336 335328
rect 287388 335316 287394 335368
rect 289078 335316 289084 335368
rect 289136 335356 289142 335368
rect 315022 335356 315028 335368
rect 289136 335328 315028 335356
rect 289136 335316 289142 335328
rect 315022 335316 315028 335328
rect 315080 335316 315086 335368
rect 316678 335316 316684 335368
rect 316736 335356 316742 335368
rect 343358 335356 343364 335368
rect 316736 335328 343364 335356
rect 316736 335316 316742 335328
rect 343358 335316 343364 335328
rect 343416 335316 343422 335368
rect 344278 335316 344284 335368
rect 344336 335356 344342 335368
rect 371326 335356 371332 335368
rect 344336 335328 371332 335356
rect 344336 335316 344342 335328
rect 371326 335316 371332 335328
rect 371384 335316 371390 335368
rect 373258 335316 373264 335368
rect 373316 335356 373322 335368
rect 399018 335356 399024 335368
rect 373316 335328 399024 335356
rect 373316 335316 373322 335328
rect 399018 335316 399024 335328
rect 399076 335316 399082 335368
rect 400858 335316 400864 335368
rect 400916 335356 400922 335368
rect 427354 335356 427360 335368
rect 400916 335328 427360 335356
rect 400916 335316 400922 335328
rect 427354 335316 427360 335328
rect 427412 335316 427418 335368
rect 428458 335316 428464 335368
rect 428516 335356 428522 335368
rect 455322 335356 455328 335368
rect 428516 335328 455328 335356
rect 428516 335316 428522 335328
rect 455322 335316 455328 335328
rect 455380 335316 455386 335368
rect 456058 335316 456064 335368
rect 456116 335356 456122 335368
rect 483198 335356 483204 335368
rect 456116 335328 483204 335356
rect 456116 335316 456122 335328
rect 483198 335316 483204 335328
rect 483256 335316 483262 335368
rect 485038 335316 485044 335368
rect 485096 335356 485102 335368
rect 511350 335356 511356 335368
rect 485096 335328 511356 335356
rect 485096 335316 485102 335328
rect 511350 335316 511356 335328
rect 511408 335316 511414 335368
rect 512638 335316 512644 335368
rect 512696 335356 512702 335368
rect 539318 335356 539324 335368
rect 512696 335328 539324 335356
rect 512696 335316 512702 335328
rect 539318 335316 539324 335328
rect 539376 335316 539382 335368
rect 540238 335316 540244 335368
rect 540296 335356 540302 335368
rect 567194 335356 567200 335368
rect 540296 335328 567200 335356
rect 540296 335316 540302 335328
rect 567194 335316 567200 335328
rect 567252 335316 567258 335368
rect 37918 333208 37924 333260
rect 37976 333248 37982 333260
rect 545758 333248 545764 333260
rect 37976 333220 545764 333248
rect 37976 333208 37982 333220
rect 545758 333208 545764 333220
rect 545816 333208 545822 333260
rect 35618 332528 35624 332580
rect 35676 332568 35682 332580
rect 36814 332568 36820 332580
rect 35676 332540 36820 332568
rect 35676 332528 35682 332540
rect 36814 332528 36820 332540
rect 36872 332528 36878 332580
rect 209682 331236 209688 331288
rect 209740 331276 209746 331288
rect 262214 331276 262220 331288
rect 209740 331248 262220 331276
rect 209740 331236 209746 331248
rect 262214 331236 262220 331248
rect 262272 331236 262278 331288
rect 266262 331236 266268 331288
rect 266320 331276 266326 331288
rect 317414 331276 317420 331288
rect 266320 331248 317420 331276
rect 266320 331236 266326 331248
rect 317414 331236 317420 331248
rect 317472 331236 317478 331288
rect 405642 331236 405648 331288
rect 405700 331276 405706 331288
rect 458174 331276 458180 331288
rect 405700 331248 458180 331276
rect 405700 331236 405706 331248
rect 458174 331236 458180 331248
rect 458232 331236 458238 331288
rect 462222 331236 462228 331288
rect 462280 331276 462286 331288
rect 513374 331276 513380 331288
rect 462280 331248 513380 331276
rect 462280 331236 462286 331248
rect 513374 331236 513380 331248
rect 513432 331236 513438 331288
rect 483658 315936 483664 315988
rect 483716 315976 483722 315988
rect 491662 315976 491668 315988
rect 483716 315948 491668 315976
rect 483716 315936 483722 315948
rect 491662 315936 491668 315948
rect 491720 315936 491726 315988
rect 428642 315256 428648 315308
rect 428700 315296 428706 315308
rect 435726 315296 435732 315308
rect 428700 315268 435732 315296
rect 428700 315256 428706 315268
rect 435726 315256 435732 315268
rect 435784 315256 435790 315308
rect 512730 315256 512736 315308
rect 512788 315296 512794 315308
rect 519630 315296 519636 315308
rect 512788 315268 519636 315296
rect 512788 315256 512794 315268
rect 519630 315256 519636 315268
rect 519688 315256 519694 315308
rect 232682 315120 232688 315172
rect 232740 315160 232746 315172
rect 239766 315160 239772 315172
rect 232740 315132 239772 315160
rect 232740 315120 232746 315132
rect 239766 315120 239772 315132
rect 239824 315120 239830 315172
rect 63586 314644 63592 314696
rect 63644 314684 63650 314696
rect 64322 314684 64328 314696
rect 63644 314656 64328 314684
rect 63644 314644 63650 314656
rect 64322 314644 64328 314656
rect 64380 314644 64386 314696
rect 287698 314644 287704 314696
rect 287756 314684 287762 314696
rect 295702 314684 295708 314696
rect 287756 314656 295708 314684
rect 287756 314644 287762 314656
rect 295702 314644 295708 314656
rect 295760 314644 295766 314696
rect 316770 314644 316776 314696
rect 316828 314684 316834 314696
rect 323670 314684 323676 314696
rect 316828 314656 323676 314684
rect 316828 314644 316834 314656
rect 323670 314644 323676 314656
rect 323728 314644 323734 314696
rect 13722 314576 13728 314628
rect 13780 314616 13786 314628
rect 66254 314616 66260 314628
rect 13780 314588 66260 314616
rect 13780 314576 13786 314588
rect 66254 314576 66260 314588
rect 66312 314576 66318 314628
rect 70302 314576 70308 314628
rect 70360 314616 70366 314628
rect 121454 314616 121460 314628
rect 70360 314588 121460 314616
rect 70360 314576 70366 314588
rect 121454 314576 121460 314588
rect 121512 314576 121518 314628
rect 126882 314576 126888 314628
rect 126940 314616 126946 314628
rect 178034 314616 178040 314628
rect 126940 314588 178040 314616
rect 126940 314576 126946 314588
rect 178034 314576 178040 314588
rect 178092 314576 178098 314628
rect 182082 314576 182088 314628
rect 182140 314616 182146 314628
rect 233234 314616 233240 314628
rect 182140 314588 233240 314616
rect 182140 314576 182146 314588
rect 233234 314576 233240 314588
rect 233292 314576 233298 314628
rect 238662 314576 238668 314628
rect 238720 314616 238726 314628
rect 289814 314616 289820 314628
rect 238720 314588 289820 314616
rect 238720 314576 238726 314588
rect 289814 314576 289820 314588
rect 289872 314576 289878 314628
rect 293862 314576 293868 314628
rect 293920 314616 293926 314628
rect 345014 314616 345020 314628
rect 293920 314588 345020 314616
rect 293920 314576 293926 314588
rect 345014 314576 345020 314588
rect 345072 314576 345078 314628
rect 350442 314576 350448 314628
rect 350500 314616 350506 314628
rect 401594 314616 401600 314628
rect 350500 314588 401600 314616
rect 350500 314576 350506 314588
rect 401594 314576 401600 314588
rect 401652 314576 401658 314628
rect 427722 314576 427728 314628
rect 427780 314616 427786 314628
rect 428550 314616 428556 314628
rect 427780 314588 428556 314616
rect 427780 314576 427786 314588
rect 428550 314576 428556 314588
rect 428608 314576 428614 314628
rect 434622 314576 434628 314628
rect 434680 314616 434686 314628
rect 485774 314616 485780 314628
rect 434680 314588 485780 314616
rect 434680 314576 434686 314588
rect 485774 314576 485780 314588
rect 485832 314576 485838 314628
rect 489822 314576 489828 314628
rect 489880 314616 489886 314628
rect 542354 314616 542360 314628
rect 489880 314588 542360 314616
rect 489880 314576 489886 314588
rect 542354 314576 542360 314588
rect 542412 314576 542418 314628
rect 35618 314508 35624 314560
rect 35676 314548 35682 314560
rect 36998 314548 37004 314560
rect 35676 314520 37004 314548
rect 35676 314508 35682 314520
rect 36998 314508 37004 314520
rect 37056 314508 37062 314560
rect 42702 314508 42708 314560
rect 42760 314548 42766 314560
rect 93854 314548 93860 314560
rect 42760 314520 93860 314548
rect 42760 314508 42766 314520
rect 93854 314508 93860 314520
rect 93912 314508 93918 314560
rect 97902 314508 97908 314560
rect 97960 314548 97966 314560
rect 149054 314548 149060 314560
rect 97960 314520 149060 314548
rect 97960 314508 97966 314520
rect 149054 314508 149060 314520
rect 149112 314508 149118 314560
rect 154482 314508 154488 314560
rect 154540 314548 154546 314560
rect 205634 314548 205640 314560
rect 154540 314520 205640 314548
rect 154540 314508 154546 314520
rect 205634 314508 205640 314520
rect 205692 314508 205698 314560
rect 259730 314508 259736 314560
rect 259788 314548 259794 314560
rect 260190 314548 260196 314560
rect 259788 314520 260196 314548
rect 259788 314508 259794 314520
rect 260190 314508 260196 314520
rect 260248 314508 260254 314560
rect 322842 314508 322848 314560
rect 322900 314548 322906 314560
rect 373994 314548 374000 314560
rect 322900 314520 374000 314548
rect 322900 314508 322906 314520
rect 373994 314508 374000 314520
rect 374052 314508 374058 314560
rect 378042 314508 378048 314560
rect 378100 314548 378106 314560
rect 429194 314548 429200 314560
rect 378100 314520 429200 314548
rect 378100 314508 378106 314520
rect 429194 314508 429200 314520
rect 429252 314508 429258 314560
rect 455690 314508 455696 314560
rect 455748 314548 455754 314560
rect 456150 314548 456156 314560
rect 455748 314520 456156 314548
rect 455748 314508 455754 314520
rect 456150 314508 456156 314520
rect 456208 314508 456214 314560
rect 518802 314508 518808 314560
rect 518860 314548 518866 314560
rect 569954 314548 569960 314560
rect 518860 314520 569960 314548
rect 518860 314508 518866 314520
rect 569954 314508 569960 314520
rect 570012 314508 570018 314560
rect 343542 314440 343548 314492
rect 343600 314480 343606 314492
rect 345658 314480 345664 314492
rect 343600 314452 345664 314480
rect 343600 314440 343606 314452
rect 345658 314440 345664 314452
rect 345716 314440 345722 314492
rect 25682 311788 25688 311840
rect 25740 311828 25746 311840
rect 36722 311828 36728 311840
rect 25740 311800 36728 311828
rect 25740 311788 25746 311800
rect 36722 311788 36728 311800
rect 36780 311788 36786 311840
rect 42886 311788 42892 311840
rect 42944 311828 42950 311840
rect 72050 311828 72056 311840
rect 42944 311800 45554 311828
rect 42944 311788 42950 311800
rect 15194 311720 15200 311772
rect 15252 311760 15258 311772
rect 43990 311760 43996 311772
rect 15252 311732 43996 311760
rect 15252 311720 15258 311732
rect 43990 311720 43996 311732
rect 44048 311720 44054 311772
rect 45526 311760 45554 311800
rect 64846 311800 72056 311828
rect 64846 311760 64874 311800
rect 72050 311788 72056 311800
rect 72108 311788 72114 311840
rect 99466 311788 99472 311840
rect 99524 311828 99530 311840
rect 99524 311800 103514 311828
rect 99524 311788 99530 311800
rect 45526 311732 64874 311760
rect 71866 311720 71872 311772
rect 71924 311760 71930 311772
rect 100018 311760 100024 311772
rect 71924 311732 100024 311760
rect 71924 311720 71930 311732
rect 100018 311720 100024 311732
rect 100076 311720 100082 311772
rect 103486 311760 103514 311800
rect 127066 311788 127072 311840
rect 127124 311828 127130 311840
rect 127124 311800 132494 311828
rect 127124 311788 127130 311800
rect 127986 311760 127992 311772
rect 103486 311732 127992 311760
rect 127986 311720 127992 311732
rect 128044 311720 128050 311772
rect 132466 311760 132494 311800
rect 183646 311788 183652 311840
rect 183704 311828 183710 311840
rect 183704 311800 190454 311828
rect 183704 311788 183710 311800
rect 156046 311760 156052 311772
rect 132466 311732 156052 311760
rect 156046 311720 156052 311732
rect 156104 311720 156110 311772
rect 165982 311720 165988 311772
rect 166040 311760 166046 311772
rect 177298 311760 177304 311772
rect 166040 311732 177304 311760
rect 166040 311720 166046 311732
rect 177298 311720 177304 311732
rect 177356 311720 177362 311772
rect 178678 311720 178684 311772
rect 178736 311760 178742 311772
rect 184014 311760 184020 311772
rect 178736 311732 184020 311760
rect 178736 311720 178742 311732
rect 184014 311720 184020 311732
rect 184072 311720 184078 311772
rect 190426 311760 190454 311800
rect 374638 311788 374644 311840
rect 374696 311828 374702 311840
rect 379698 311828 379704 311840
rect 374696 311800 379704 311828
rect 374696 311788 374702 311800
rect 379698 311788 379704 311800
rect 379756 311788 379762 311840
rect 539318 311788 539324 311840
rect 539376 311828 539382 311840
rect 542998 311828 543004 311840
rect 539376 311800 543004 311828
rect 539376 311788 539382 311800
rect 542998 311788 543004 311800
rect 543056 311788 543062 311840
rect 211706 311760 211712 311772
rect 190426 311732 211712 311760
rect 211706 311720 211712 311732
rect 211764 311720 211770 311772
rect 222010 311720 222016 311772
rect 222068 311760 222074 311772
rect 232590 311760 232596 311772
rect 222068 311732 232596 311760
rect 222068 311720 222074 311732
rect 232590 311720 232596 311732
rect 232648 311720 232654 311772
rect 249702 311720 249708 311772
rect 249760 311760 249766 311772
rect 260098 311760 260104 311772
rect 249760 311732 260104 311760
rect 249760 311720 249766 311732
rect 260098 311720 260104 311732
rect 260156 311720 260162 311772
rect 261478 311720 261484 311772
rect 261536 311760 261542 311772
rect 567194 311760 567200 311772
rect 261536 311732 567200 311760
rect 261536 311720 261542 311732
rect 567194 311720 567200 311732
rect 567252 311720 567258 311772
rect 53650 311652 53656 311704
rect 53708 311692 53714 311704
rect 69658 311692 69664 311704
rect 53708 311664 69664 311692
rect 53708 311652 53714 311664
rect 69658 311652 69664 311664
rect 69716 311652 69722 311704
rect 81986 311652 81992 311704
rect 82044 311692 82050 311704
rect 94498 311692 94504 311704
rect 82044 311664 94504 311692
rect 82044 311652 82050 311664
rect 94498 311652 94504 311664
rect 94556 311652 94562 311704
rect 109678 311652 109684 311704
rect 109736 311692 109742 311704
rect 120718 311692 120724 311704
rect 109736 311664 120724 311692
rect 109736 311652 109742 311664
rect 120718 311652 120724 311664
rect 120776 311652 120782 311704
rect 137646 311652 137652 311704
rect 137704 311692 137710 311704
rect 148410 311692 148416 311704
rect 137704 311664 148416 311692
rect 137704 311652 137710 311664
rect 148410 311652 148416 311664
rect 148468 311652 148474 311704
rect 193674 311652 193680 311704
rect 193732 311692 193738 311704
rect 204898 311692 204904 311704
rect 193732 311664 204904 311692
rect 193732 311652 193738 311664
rect 204898 311652 204904 311664
rect 204956 311652 204962 311704
rect 238846 311652 238852 311704
rect 238904 311692 238910 311704
rect 268010 311692 268016 311704
rect 238904 311664 268016 311692
rect 238904 311652 238910 311664
rect 268010 311652 268016 311664
rect 268068 311652 268074 311704
rect 277670 311652 277676 311704
rect 277728 311692 277734 311704
rect 289078 311692 289084 311704
rect 277728 311664 289084 311692
rect 277728 311652 277734 311664
rect 289078 311652 289084 311664
rect 289136 311652 289142 311704
rect 306006 311652 306012 311704
rect 306064 311692 306070 311704
rect 316678 311692 316684 311704
rect 306064 311664 316684 311692
rect 306064 311652 306070 311664
rect 316678 311652 316684 311664
rect 316736 311652 316742 311704
rect 323026 311652 323032 311704
rect 323084 311692 323090 311704
rect 352006 311692 352012 311704
rect 323084 311664 352012 311692
rect 323084 311652 323090 311664
rect 352006 311652 352012 311664
rect 352064 311652 352070 311704
rect 361666 311652 361672 311704
rect 361724 311692 361730 311704
rect 373258 311692 373264 311704
rect 361724 311664 373264 311692
rect 361724 311652 361730 311664
rect 373258 311652 373264 311664
rect 373316 311652 373322 311704
rect 379606 311652 379612 311704
rect 379664 311692 379670 311704
rect 408034 311692 408040 311704
rect 379664 311664 408040 311692
rect 379664 311652 379670 311664
rect 408034 311652 408040 311664
rect 408092 311652 408098 311704
rect 417694 311652 417700 311704
rect 417752 311692 417758 311704
rect 428458 311692 428464 311704
rect 417752 311664 428464 311692
rect 417752 311652 417758 311664
rect 428458 311652 428464 311664
rect 428516 311652 428522 311704
rect 434806 311652 434812 311704
rect 434864 311692 434870 311704
rect 463694 311692 463700 311704
rect 434864 311664 463700 311692
rect 434864 311652 434870 311664
rect 463694 311652 463700 311664
rect 463752 311652 463758 311704
rect 473998 311652 474004 311704
rect 474056 311692 474062 311704
rect 485038 311692 485044 311704
rect 474056 311664 485044 311692
rect 474056 311652 474062 311664
rect 485038 311652 485044 311664
rect 485096 311652 485102 311704
rect 501690 311652 501696 311704
rect 501748 311692 501754 311704
rect 512638 311692 512644 311704
rect 501748 311664 512644 311692
rect 501748 311652 501754 311664
rect 512638 311652 512644 311664
rect 512696 311652 512702 311704
rect 518986 311652 518992 311704
rect 519044 311692 519050 311704
rect 547874 311692 547880 311704
rect 519044 311664 547880 311692
rect 519044 311652 519050 311664
rect 547874 311652 547880 311664
rect 547932 311652 547938 311704
rect 333698 311584 333704 311636
rect 333756 311624 333762 311636
rect 344278 311624 344284 311636
rect 333756 311596 344284 311624
rect 333756 311584 333762 311596
rect 344278 311584 344284 311596
rect 344336 311584 344342 311636
rect 390002 311584 390008 311636
rect 390060 311624 390066 311636
rect 400858 311624 400864 311636
rect 390060 311596 400864 311624
rect 390060 311584 390066 311596
rect 400858 311584 400864 311596
rect 400916 311584 400922 311636
rect 445662 311584 445668 311636
rect 445720 311624 445726 311636
rect 456058 311624 456064 311636
rect 445720 311596 456064 311624
rect 445720 311584 445726 311596
rect 456058 311584 456064 311596
rect 456116 311584 456122 311636
rect 529658 311584 529664 311636
rect 529716 311624 529722 311636
rect 540238 311624 540244 311636
rect 529716 311596 540244 311624
rect 529716 311584 529722 311596
rect 540238 311584 540244 311596
rect 540296 311584 540302 311636
rect 36906 311516 36912 311568
rect 36964 311556 36970 311568
rect 557534 311556 557540 311568
rect 36964 311528 557540 311556
rect 36964 311516 36970 311528
rect 557534 311516 557540 311528
rect 557592 311516 557598 311568
rect 16022 308388 16028 308440
rect 16080 308428 16086 308440
rect 547874 308428 547880 308440
rect 16080 308400 547880 308428
rect 16080 308388 16086 308400
rect 547874 308388 547880 308400
rect 547932 308388 547938 308440
rect 25682 308048 25688 308100
rect 25740 308088 25746 308100
rect 261478 308088 261484 308100
rect 25740 308060 261484 308088
rect 25740 308048 25746 308060
rect 261478 308048 261484 308060
rect 261536 308048 261542 308100
rect 148318 307980 148324 308032
rect 148376 308020 148382 308032
rect 165614 308020 165620 308032
rect 148376 307992 165620 308020
rect 148376 307980 148382 307992
rect 165614 307980 165620 307992
rect 165672 307980 165678 308032
rect 175458 307980 175464 308032
rect 175516 308020 175522 308032
rect 193674 308020 193680 308032
rect 175516 307992 193680 308020
rect 175516 307980 175522 307992
rect 193674 307980 193680 307992
rect 193732 307980 193738 308032
rect 203518 307980 203524 308032
rect 203576 308020 203582 308032
rect 221366 308020 221372 308032
rect 203576 307992 221372 308020
rect 203576 307980 203582 307992
rect 221366 307980 221372 307992
rect 221424 307980 221430 308032
rect 296346 307980 296352 308032
rect 296404 308020 296410 308032
rect 316770 308020 316776 308032
rect 296404 307992 316776 308020
rect 296404 307980 296410 307992
rect 316770 307980 316776 307992
rect 316828 307980 316834 308032
rect 408034 307980 408040 308032
rect 408092 308020 408098 308032
rect 428642 308020 428648 308032
rect 408092 307992 428648 308020
rect 408092 307980 408098 307992
rect 428642 307980 428648 307992
rect 428700 307980 428706 308032
rect 492030 307980 492036 308032
rect 492088 308020 492094 308032
rect 512730 308020 512736 308032
rect 492088 307992 512736 308020
rect 492088 307980 492094 307992
rect 512730 307980 512736 307992
rect 512788 307980 512794 308032
rect 36998 307912 37004 307964
rect 37056 307952 37062 307964
rect 53650 307952 53656 307964
rect 37056 307924 53656 307952
rect 37056 307912 37062 307924
rect 53650 307912 53656 307924
rect 53708 307912 53714 307964
rect 64322 307912 64328 307964
rect 64380 307952 64386 307964
rect 81434 307952 81440 307964
rect 64380 307924 81440 307952
rect 64380 307912 64386 307924
rect 81434 307912 81440 307924
rect 81492 307912 81498 307964
rect 91462 307912 91468 307964
rect 91520 307952 91526 307964
rect 109678 307952 109684 307964
rect 91520 307924 109684 307952
rect 91520 307912 91526 307924
rect 109678 307912 109684 307924
rect 109736 307912 109742 307964
rect 119430 307912 119436 307964
rect 119488 307952 119494 307964
rect 137646 307952 137652 307964
rect 119488 307924 137652 307952
rect 119488 307912 119494 307924
rect 137646 307912 137652 307924
rect 137704 307912 137710 307964
rect 156322 307912 156328 307964
rect 156380 307952 156386 307964
rect 178678 307952 178684 307964
rect 156380 307924 178684 307952
rect 156380 307912 156386 307924
rect 178678 307912 178684 307924
rect 178736 307912 178742 307964
rect 232590 307912 232596 307964
rect 232648 307952 232654 307964
rect 249702 307952 249708 307964
rect 232648 307924 249708 307952
rect 232648 307912 232654 307924
rect 249702 307912 249708 307924
rect 249760 307912 249766 307964
rect 260190 307912 260196 307964
rect 260248 307952 260254 307964
rect 277670 307952 277676 307964
rect 260248 307924 277676 307952
rect 260248 307912 260254 307924
rect 277670 307912 277676 307924
rect 277728 307912 277734 307964
rect 287514 307912 287520 307964
rect 287572 307952 287578 307964
rect 305362 307952 305368 307964
rect 287572 307924 305368 307952
rect 287572 307912 287578 307924
rect 305362 307912 305368 307924
rect 305420 307912 305426 307964
rect 345658 307912 345664 307964
rect 345716 307952 345722 307964
rect 361666 307952 361672 307964
rect 345716 307924 361672 307952
rect 345716 307912 345722 307924
rect 361666 307912 361672 307924
rect 361724 307912 361730 307964
rect 371510 307912 371516 307964
rect 371568 307952 371574 307964
rect 389358 307952 389364 307964
rect 371568 307924 389364 307952
rect 371568 307912 371574 307924
rect 389358 307912 389364 307924
rect 389416 307912 389422 307964
rect 399478 307912 399484 307964
rect 399536 307952 399542 307964
rect 417694 307952 417700 307964
rect 399536 307924 417700 307952
rect 399536 307912 399542 307924
rect 417694 307912 417700 307924
rect 417752 307912 417758 307964
rect 456058 307912 456064 307964
rect 456116 307952 456122 307964
rect 473538 307952 473544 307964
rect 456116 307924 473544 307952
rect 456116 307912 456122 307924
rect 473538 307912 473544 307924
rect 473596 307912 473602 307964
rect 483474 307912 483480 307964
rect 483532 307952 483538 307964
rect 501690 307952 501696 307964
rect 483532 307924 501696 307952
rect 483532 307912 483538 307924
rect 501690 307912 501696 307924
rect 501748 307912 501754 307964
rect 36906 307844 36912 307896
rect 36964 307884 36970 307896
rect 63310 307884 63316 307896
rect 36964 307856 63316 307884
rect 36964 307844 36970 307856
rect 63310 307844 63316 307856
rect 63368 307844 63374 307896
rect 66898 307844 66904 307896
rect 66956 307884 66962 307896
rect 91094 307884 91100 307896
rect 66956 307856 91100 307884
rect 66956 307844 66962 307856
rect 91094 307844 91100 307856
rect 91152 307844 91158 307896
rect 94498 307844 94504 307896
rect 94556 307884 94562 307896
rect 119338 307884 119344 307896
rect 94556 307856 119344 307884
rect 94556 307844 94562 307856
rect 119338 307844 119344 307856
rect 119396 307844 119402 307896
rect 120718 307844 120724 307896
rect 120776 307884 120782 307896
rect 147306 307884 147312 307896
rect 120776 307856 147312 307884
rect 120776 307844 120782 307856
rect 147306 307844 147312 307856
rect 147364 307844 147370 307896
rect 148410 307844 148416 307896
rect 148468 307884 148474 307896
rect 175274 307884 175280 307896
rect 148468 307856 175280 307884
rect 148468 307844 148474 307856
rect 175274 307844 175280 307856
rect 175332 307844 175338 307896
rect 177298 307844 177304 307896
rect 177356 307884 177362 307896
rect 203334 307884 203340 307896
rect 177356 307856 203340 307884
rect 177356 307844 177362 307856
rect 203334 307844 203340 307856
rect 203392 307844 203398 307896
rect 204898 307844 204904 307896
rect 204956 307884 204962 307896
rect 231026 307884 231032 307896
rect 204956 307856 231032 307884
rect 204956 307844 204962 307856
rect 231026 307844 231032 307856
rect 231084 307844 231090 307896
rect 232498 307844 232504 307896
rect 232556 307884 232562 307896
rect 259362 307884 259368 307896
rect 232556 307856 259368 307884
rect 232556 307844 232562 307856
rect 259362 307844 259368 307856
rect 259420 307844 259426 307896
rect 268010 307844 268016 307896
rect 268068 307884 268074 307896
rect 287698 307884 287704 307896
rect 268068 307856 287704 307884
rect 268068 307844 268074 307856
rect 287698 307844 287704 307856
rect 287756 307844 287762 307896
rect 315482 307844 315488 307896
rect 315540 307884 315546 307896
rect 333698 307884 333704 307896
rect 315540 307856 333704 307884
rect 315540 307844 315546 307856
rect 333698 307844 333704 307856
rect 333756 307844 333762 307896
rect 352006 307844 352012 307896
rect 352064 307884 352070 307896
rect 374638 307884 374644 307896
rect 352064 307856 374644 307884
rect 352064 307844 352070 307856
rect 374638 307844 374644 307856
rect 374696 307844 374702 307896
rect 428550 307844 428556 307896
rect 428608 307884 428614 307896
rect 445662 307884 445668 307896
rect 428608 307856 445668 307884
rect 428608 307844 428614 307856
rect 445662 307844 445668 307856
rect 445720 307844 445726 307896
rect 464338 307844 464344 307896
rect 464396 307884 464402 307896
rect 483658 307884 483664 307896
rect 464396 307856 483664 307884
rect 464396 307844 464402 307856
rect 483658 307844 483664 307856
rect 483716 307844 483722 307896
rect 511442 307844 511448 307896
rect 511500 307884 511506 307896
rect 529658 307884 529664 307896
rect 511500 307856 529664 307884
rect 511500 307844 511506 307856
rect 529658 307844 529664 307856
rect 529716 307844 529722 307896
rect 542998 307844 543004 307896
rect 543056 307884 543062 307896
rect 557534 307884 557540 307896
rect 543056 307856 557540 307884
rect 543056 307844 543062 307856
rect 557534 307844 557540 307856
rect 557592 307844 557598 307896
rect 212258 307776 212264 307828
rect 212316 307816 212322 307828
rect 232682 307816 232688 307828
rect 212316 307788 232688 307816
rect 212316 307776 212322 307788
rect 232682 307776 232688 307788
rect 232740 307776 232746 307828
rect 260098 307776 260104 307828
rect 260156 307816 260162 307828
rect 287330 307816 287336 307828
rect 260156 307788 287336 307816
rect 260156 307776 260162 307788
rect 287330 307776 287336 307788
rect 287388 307776 287394 307828
rect 289078 307776 289084 307828
rect 289136 307816 289142 307828
rect 315022 307816 315028 307828
rect 289136 307788 315028 307816
rect 289136 307776 289142 307788
rect 315022 307776 315028 307788
rect 315080 307776 315086 307828
rect 316678 307776 316684 307828
rect 316736 307816 316742 307828
rect 343358 307816 343364 307828
rect 316736 307788 343364 307816
rect 316736 307776 316742 307788
rect 343358 307776 343364 307788
rect 343416 307776 343422 307828
rect 344278 307776 344284 307828
rect 344336 307816 344342 307828
rect 371326 307816 371332 307828
rect 344336 307788 371332 307816
rect 344336 307776 344342 307788
rect 371326 307776 371332 307788
rect 371384 307776 371390 307828
rect 373258 307776 373264 307828
rect 373316 307816 373322 307828
rect 399018 307816 399024 307828
rect 373316 307788 399024 307816
rect 373316 307776 373322 307788
rect 399018 307776 399024 307788
rect 399076 307776 399082 307828
rect 400858 307776 400864 307828
rect 400916 307816 400922 307828
rect 427354 307816 427360 307828
rect 400916 307788 427360 307816
rect 400916 307776 400922 307788
rect 427354 307776 427360 307788
rect 427412 307776 427418 307828
rect 428458 307776 428464 307828
rect 428516 307816 428522 307828
rect 455322 307816 455328 307828
rect 428516 307788 455328 307816
rect 428516 307776 428522 307788
rect 455322 307776 455328 307788
rect 455380 307776 455386 307828
rect 456150 307776 456156 307828
rect 456208 307816 456214 307828
rect 483198 307816 483204 307828
rect 456208 307788 483204 307816
rect 456208 307776 456214 307788
rect 483198 307776 483204 307788
rect 483256 307776 483262 307828
rect 485038 307776 485044 307828
rect 485096 307816 485102 307828
rect 511350 307816 511356 307828
rect 485096 307788 511356 307816
rect 485096 307776 485102 307788
rect 511350 307776 511356 307788
rect 511408 307776 511414 307828
rect 512638 307776 512644 307828
rect 512696 307816 512702 307828
rect 539318 307816 539324 307828
rect 512696 307788 539324 307816
rect 512696 307776 512702 307788
rect 539318 307776 539324 307788
rect 539376 307776 539382 307828
rect 540238 307776 540244 307828
rect 540296 307816 540302 307828
rect 567194 307816 567200 307828
rect 540296 307788 567200 307816
rect 540296 307776 540302 307788
rect 567194 307776 567200 307788
rect 567252 307776 567258 307828
rect 37918 305600 37924 305652
rect 37976 305640 37982 305652
rect 545758 305640 545764 305652
rect 37976 305612 545764 305640
rect 37976 305600 37982 305612
rect 545758 305600 545764 305612
rect 545816 305600 545822 305652
rect 3050 304988 3056 305040
rect 3108 305028 3114 305040
rect 10318 305028 10324 305040
rect 3108 305000 10324 305028
rect 3108 304988 3114 305000
rect 10318 304988 10324 305000
rect 10376 304988 10382 305040
rect 35618 304988 35624 305040
rect 35676 305028 35682 305040
rect 36722 305028 36728 305040
rect 35676 305000 36728 305028
rect 35676 304988 35682 305000
rect 36722 304988 36728 305000
rect 36780 304988 36786 305040
rect 63586 291864 63592 291916
rect 63644 291904 63650 291916
rect 64322 291904 64328 291916
rect 63644 291876 64328 291904
rect 63644 291864 63650 291876
rect 64322 291864 64328 291876
rect 64380 291864 64386 291916
rect 259730 291864 259736 291916
rect 259788 291904 259794 291916
rect 260190 291904 260196 291916
rect 259788 291876 260196 291904
rect 259788 291864 259794 291876
rect 260190 291864 260196 291876
rect 260248 291864 260254 291916
rect 287698 288328 287704 288380
rect 287756 288368 287762 288380
rect 295702 288368 295708 288380
rect 287756 288340 295708 288368
rect 287756 288328 287762 288340
rect 295702 288328 295708 288340
rect 295760 288328 295766 288380
rect 316770 288328 316776 288380
rect 316828 288368 316834 288380
rect 323670 288368 323676 288380
rect 316828 288340 323676 288368
rect 316828 288328 316834 288340
rect 323670 288328 323676 288340
rect 323728 288328 323734 288380
rect 232682 287920 232688 287972
rect 232740 287960 232746 287972
rect 239766 287960 239772 287972
rect 232740 287932 239772 287960
rect 232740 287920 232746 287932
rect 239766 287920 239772 287932
rect 239824 287920 239830 287972
rect 428642 287648 428648 287700
rect 428700 287688 428706 287700
rect 435726 287688 435732 287700
rect 428700 287660 435732 287688
rect 428700 287648 428706 287660
rect 435726 287648 435732 287660
rect 435784 287648 435790 287700
rect 512730 287512 512736 287564
rect 512788 287552 512794 287564
rect 519630 287552 519636 287564
rect 512788 287524 519636 287552
rect 512788 287512 512794 287524
rect 519630 287512 519636 287524
rect 519688 287512 519694 287564
rect 483658 287376 483664 287428
rect 483716 287416 483722 287428
rect 491662 287416 491668 287428
rect 483716 287388 491668 287416
rect 483716 287376 483722 287388
rect 491662 287376 491668 287388
rect 491720 287376 491726 287428
rect 13722 286968 13728 287020
rect 13780 287008 13786 287020
rect 66254 287008 66260 287020
rect 13780 286980 66260 287008
rect 13780 286968 13786 286980
rect 66254 286968 66260 286980
rect 66312 286968 66318 287020
rect 70302 286968 70308 287020
rect 70360 287008 70366 287020
rect 121454 287008 121460 287020
rect 70360 286980 121460 287008
rect 70360 286968 70366 286980
rect 121454 286968 121460 286980
rect 121512 286968 121518 287020
rect 126882 286968 126888 287020
rect 126940 287008 126946 287020
rect 178034 287008 178040 287020
rect 126940 286980 178040 287008
rect 126940 286968 126946 286980
rect 178034 286968 178040 286980
rect 178092 286968 178098 287020
rect 209682 286968 209688 287020
rect 209740 287008 209746 287020
rect 262214 287008 262220 287020
rect 209740 286980 262220 287008
rect 209740 286968 209746 286980
rect 262214 286968 262220 286980
rect 262272 286968 262278 287020
rect 266262 286968 266268 287020
rect 266320 287008 266326 287020
rect 317414 287008 317420 287020
rect 266320 286980 317420 287008
rect 266320 286968 266326 286980
rect 317414 286968 317420 286980
rect 317472 286968 317478 287020
rect 322842 286968 322848 287020
rect 322900 287008 322906 287020
rect 373994 287008 374000 287020
rect 322900 286980 374000 287008
rect 322900 286968 322906 286980
rect 373994 286968 374000 286980
rect 374052 286968 374058 287020
rect 405642 286968 405648 287020
rect 405700 287008 405706 287020
rect 458174 287008 458180 287020
rect 405700 286980 458180 287008
rect 405700 286968 405706 286980
rect 458174 286968 458180 286980
rect 458232 286968 458238 287020
rect 489822 286968 489828 287020
rect 489880 287008 489886 287020
rect 542354 287008 542360 287020
rect 489880 286980 542360 287008
rect 489880 286968 489886 286980
rect 542354 286968 542360 286980
rect 542412 286968 542418 287020
rect 35618 286900 35624 286952
rect 35676 286940 35682 286952
rect 36998 286940 37004 286952
rect 35676 286912 37004 286940
rect 35676 286900 35682 286912
rect 36998 286900 37004 286912
rect 37056 286900 37062 286952
rect 42702 286900 42708 286952
rect 42760 286940 42766 286952
rect 93854 286940 93860 286952
rect 42760 286912 93860 286940
rect 42760 286900 42766 286912
rect 93854 286900 93860 286912
rect 93912 286900 93918 286952
rect 97902 286900 97908 286952
rect 97960 286940 97966 286952
rect 149054 286940 149060 286952
rect 97960 286912 149060 286940
rect 97960 286900 97966 286912
rect 149054 286900 149060 286912
rect 149112 286900 149118 286952
rect 154482 286900 154488 286952
rect 154540 286940 154546 286952
rect 205634 286940 205640 286952
rect 154540 286912 205640 286940
rect 154540 286900 154546 286912
rect 205634 286900 205640 286912
rect 205692 286900 205698 286952
rect 238662 286900 238668 286952
rect 238720 286940 238726 286952
rect 289814 286940 289820 286952
rect 238720 286912 289820 286940
rect 238720 286900 238726 286912
rect 289814 286900 289820 286912
rect 289872 286900 289878 286952
rect 293862 286900 293868 286952
rect 293920 286940 293926 286952
rect 293920 286912 335354 286940
rect 293920 286900 293926 286912
rect 182082 286832 182088 286884
rect 182140 286872 182146 286884
rect 233234 286872 233240 286884
rect 182140 286844 233240 286872
rect 182140 286832 182146 286844
rect 233234 286832 233240 286844
rect 233292 286832 233298 286884
rect 335326 286872 335354 286912
rect 343542 286900 343548 286952
rect 343600 286940 343606 286952
rect 345658 286940 345664 286952
rect 343600 286912 345664 286940
rect 343600 286900 343606 286912
rect 345658 286900 345664 286912
rect 345716 286900 345722 286952
rect 350442 286900 350448 286952
rect 350500 286940 350506 286952
rect 401594 286940 401600 286952
rect 350500 286912 401600 286940
rect 350500 286900 350506 286912
rect 401594 286900 401600 286912
rect 401652 286900 401658 286952
rect 434622 286900 434628 286952
rect 434680 286940 434686 286952
rect 485774 286940 485780 286952
rect 434680 286912 485780 286940
rect 434680 286900 434686 286912
rect 485774 286900 485780 286912
rect 485832 286900 485838 286952
rect 518802 286900 518808 286952
rect 518860 286940 518866 286952
rect 569954 286940 569960 286952
rect 518860 286912 569960 286940
rect 518860 286900 518866 286912
rect 569954 286900 569960 286912
rect 570012 286900 570018 286952
rect 345014 286872 345020 286884
rect 335326 286844 345020 286872
rect 345014 286832 345020 286844
rect 345072 286832 345078 286884
rect 378042 286832 378048 286884
rect 378100 286872 378106 286884
rect 429194 286872 429200 286884
rect 378100 286844 429200 286872
rect 378100 286832 378106 286844
rect 429194 286832 429200 286844
rect 429252 286832 429258 286884
rect 462222 286832 462228 286884
rect 462280 286872 462286 286884
rect 513374 286872 513380 286884
rect 462280 286844 513380 286872
rect 462280 286832 462286 286844
rect 513374 286832 513380 286844
rect 513432 286832 513438 286884
rect 231670 286764 231676 286816
rect 231728 286804 231734 286816
rect 232590 286804 232596 286816
rect 231728 286776 232596 286804
rect 231728 286764 231734 286776
rect 232590 286764 232596 286776
rect 232648 286764 232654 286816
rect 427722 286764 427728 286816
rect 427780 286804 427786 286816
rect 428550 286804 428556 286816
rect 427780 286776 428556 286804
rect 427780 286764 427786 286776
rect 428550 286764 428556 286776
rect 428608 286764 428614 286816
rect 539502 286764 539508 286816
rect 539560 286804 539566 286816
rect 542998 286804 543004 286816
rect 539560 286776 543004 286804
rect 539560 286764 539566 286776
rect 542998 286764 543004 286776
rect 543056 286764 543062 286816
rect 25682 284248 25688 284300
rect 25740 284288 25746 284300
rect 36906 284288 36912 284300
rect 25740 284260 36912 284288
rect 25740 284248 25746 284260
rect 36906 284248 36912 284260
rect 36964 284248 36970 284300
rect 178678 284248 178684 284300
rect 178736 284288 178742 284300
rect 184014 284288 184020 284300
rect 178736 284260 184020 284288
rect 178736 284248 178742 284260
rect 184014 284248 184020 284260
rect 184072 284248 184078 284300
rect 374638 284248 374644 284300
rect 374696 284288 374702 284300
rect 379698 284288 379704 284300
rect 374696 284260 379704 284288
rect 374696 284248 374702 284260
rect 379698 284248 379704 284260
rect 379756 284248 379762 284300
rect 15194 284180 15200 284232
rect 15252 284220 15258 284232
rect 43990 284220 43996 284232
rect 15252 284192 43996 284220
rect 15252 284180 15258 284192
rect 43990 284180 43996 284192
rect 44048 284180 44054 284232
rect 71038 284180 71044 284232
rect 71096 284220 71102 284232
rect 567194 284220 567200 284232
rect 71096 284192 567200 284220
rect 71096 284180 71102 284192
rect 567194 284180 567200 284192
rect 567252 284180 567258 284232
rect 53650 284112 53656 284164
rect 53708 284152 53714 284164
rect 66898 284152 66904 284164
rect 53708 284124 66904 284152
rect 53708 284112 53714 284124
rect 66898 284112 66904 284124
rect 66956 284112 66962 284164
rect 71866 284112 71872 284164
rect 71924 284152 71930 284164
rect 100018 284152 100024 284164
rect 71924 284124 100024 284152
rect 71924 284112 71930 284124
rect 100018 284112 100024 284124
rect 100076 284112 100082 284164
rect 127986 284152 127992 284164
rect 103486 284124 127992 284152
rect 42886 284044 42892 284096
rect 42944 284084 42950 284096
rect 72050 284084 72056 284096
rect 42944 284056 72056 284084
rect 42944 284044 42950 284056
rect 72050 284044 72056 284056
rect 72108 284044 72114 284096
rect 81986 284044 81992 284096
rect 82044 284084 82050 284096
rect 94498 284084 94504 284096
rect 82044 284056 94504 284084
rect 82044 284044 82050 284056
rect 94498 284044 94504 284056
rect 94556 284044 94562 284096
rect 99466 284044 99472 284096
rect 99524 284084 99530 284096
rect 103486 284084 103514 284124
rect 127986 284112 127992 284124
rect 128044 284112 128050 284164
rect 156046 284152 156052 284164
rect 132466 284124 156052 284152
rect 99524 284056 103514 284084
rect 99524 284044 99530 284056
rect 109678 284044 109684 284096
rect 109736 284084 109742 284096
rect 120718 284084 120724 284096
rect 109736 284056 120724 284084
rect 109736 284044 109742 284056
rect 120718 284044 120724 284056
rect 120776 284044 120782 284096
rect 127066 284044 127072 284096
rect 127124 284084 127130 284096
rect 132466 284084 132494 284124
rect 156046 284112 156052 284124
rect 156104 284112 156110 284164
rect 165982 284112 165988 284164
rect 166040 284152 166046 284164
rect 177298 284152 177304 284164
rect 166040 284124 177304 284152
rect 166040 284112 166046 284124
rect 177298 284112 177304 284124
rect 177356 284112 177362 284164
rect 183646 284112 183652 284164
rect 183704 284152 183710 284164
rect 211706 284152 211712 284164
rect 183704 284124 211712 284152
rect 183704 284112 183710 284124
rect 211706 284112 211712 284124
rect 211764 284112 211770 284164
rect 222010 284112 222016 284164
rect 222068 284152 222074 284164
rect 232498 284152 232504 284164
rect 222068 284124 232504 284152
rect 222068 284112 222074 284124
rect 232498 284112 232504 284124
rect 232556 284112 232562 284164
rect 238846 284112 238852 284164
rect 238904 284152 238910 284164
rect 268010 284152 268016 284164
rect 238904 284124 268016 284152
rect 238904 284112 238910 284124
rect 268010 284112 268016 284124
rect 268068 284112 268074 284164
rect 277670 284112 277676 284164
rect 277728 284152 277734 284164
rect 289078 284152 289084 284164
rect 277728 284124 289084 284152
rect 277728 284112 277734 284124
rect 289078 284112 289084 284124
rect 289136 284112 289142 284164
rect 306006 284112 306012 284164
rect 306064 284152 306070 284164
rect 316678 284152 316684 284164
rect 306064 284124 316684 284152
rect 306064 284112 306070 284124
rect 316678 284112 316684 284124
rect 316736 284112 316742 284164
rect 323026 284112 323032 284164
rect 323084 284152 323090 284164
rect 352006 284152 352012 284164
rect 323084 284124 352012 284152
rect 323084 284112 323090 284124
rect 352006 284112 352012 284124
rect 352064 284112 352070 284164
rect 361666 284112 361672 284164
rect 361724 284152 361730 284164
rect 373258 284152 373264 284164
rect 361724 284124 373264 284152
rect 361724 284112 361730 284124
rect 373258 284112 373264 284124
rect 373316 284112 373322 284164
rect 379606 284112 379612 284164
rect 379664 284152 379670 284164
rect 408034 284152 408040 284164
rect 379664 284124 408040 284152
rect 379664 284112 379670 284124
rect 408034 284112 408040 284124
rect 408092 284112 408098 284164
rect 417694 284112 417700 284164
rect 417752 284152 417758 284164
rect 428458 284152 428464 284164
rect 417752 284124 428464 284152
rect 417752 284112 417758 284124
rect 428458 284112 428464 284124
rect 428516 284112 428522 284164
rect 434806 284112 434812 284164
rect 434864 284152 434870 284164
rect 463694 284152 463700 284164
rect 434864 284124 463700 284152
rect 434864 284112 434870 284124
rect 463694 284112 463700 284124
rect 463752 284112 463758 284164
rect 473998 284112 474004 284164
rect 474056 284152 474062 284164
rect 485038 284152 485044 284164
rect 474056 284124 485044 284152
rect 474056 284112 474062 284124
rect 485038 284112 485044 284124
rect 485096 284112 485102 284164
rect 501690 284112 501696 284164
rect 501748 284152 501754 284164
rect 512638 284152 512644 284164
rect 501748 284124 512644 284152
rect 501748 284112 501754 284124
rect 512638 284112 512644 284124
rect 512696 284112 512702 284164
rect 518986 284112 518992 284164
rect 519044 284152 519050 284164
rect 547874 284152 547880 284164
rect 519044 284124 547880 284152
rect 519044 284112 519050 284124
rect 547874 284112 547880 284124
rect 547932 284112 547938 284164
rect 127124 284056 132494 284084
rect 127124 284044 127130 284056
rect 137646 284044 137652 284096
rect 137704 284084 137710 284096
rect 148410 284084 148416 284096
rect 137704 284056 148416 284084
rect 137704 284044 137710 284056
rect 148410 284044 148416 284056
rect 148468 284044 148474 284096
rect 193674 284044 193680 284096
rect 193732 284084 193738 284096
rect 204898 284084 204904 284096
rect 193732 284056 204904 284084
rect 193732 284044 193738 284056
rect 204898 284044 204904 284056
rect 204956 284044 204962 284096
rect 249702 284044 249708 284096
rect 249760 284084 249766 284096
rect 260098 284084 260104 284096
rect 249760 284056 260104 284084
rect 249760 284044 249766 284056
rect 260098 284044 260104 284056
rect 260156 284044 260162 284096
rect 333698 284044 333704 284096
rect 333756 284084 333762 284096
rect 344278 284084 344284 284096
rect 333756 284056 344284 284084
rect 333756 284044 333762 284056
rect 344278 284044 344284 284056
rect 344336 284044 344342 284096
rect 390002 284044 390008 284096
rect 390060 284084 390066 284096
rect 400858 284084 400864 284096
rect 390060 284056 400864 284084
rect 390060 284044 390066 284056
rect 400858 284044 400864 284056
rect 400916 284044 400922 284096
rect 445662 284044 445668 284096
rect 445720 284084 445726 284096
rect 456150 284084 456156 284096
rect 445720 284056 456156 284084
rect 445720 284044 445726 284056
rect 456150 284044 456156 284056
rect 456208 284044 456214 284096
rect 529658 284044 529664 284096
rect 529716 284084 529722 284096
rect 540238 284084 540244 284096
rect 529716 284056 540244 284084
rect 529716 284044 529722 284056
rect 540238 284044 540244 284056
rect 540296 284044 540302 284096
rect 36814 283976 36820 284028
rect 36872 284016 36878 284028
rect 557534 284016 557540 284028
rect 36872 283988 557540 284016
rect 36872 283976 36878 283988
rect 557534 283976 557540 283988
rect 557592 283976 557598 284028
rect 16022 280780 16028 280832
rect 16080 280820 16086 280832
rect 547874 280820 547880 280832
rect 16080 280792 547880 280820
rect 16080 280780 16086 280792
rect 547874 280780 547880 280792
rect 547932 280780 547938 280832
rect 25682 280372 25688 280424
rect 25740 280412 25746 280424
rect 71038 280412 71044 280424
rect 25740 280384 71044 280412
rect 25740 280372 25746 280384
rect 71038 280372 71044 280384
rect 71096 280372 71102 280424
rect 212350 280372 212356 280424
rect 212408 280412 212414 280424
rect 232682 280412 232688 280424
rect 212408 280384 232688 280412
rect 212408 280372 212414 280384
rect 232682 280372 232688 280384
rect 232740 280372 232746 280424
rect 296346 280372 296352 280424
rect 296404 280412 296410 280424
rect 316770 280412 316776 280424
rect 296404 280384 316776 280412
rect 296404 280372 296410 280384
rect 316770 280372 316776 280384
rect 316828 280372 316834 280424
rect 408034 280372 408040 280424
rect 408092 280412 408098 280424
rect 428642 280412 428648 280424
rect 408092 280384 428648 280412
rect 408092 280372 408098 280384
rect 428642 280372 428648 280384
rect 428700 280372 428706 280424
rect 492030 280372 492036 280424
rect 492088 280412 492094 280424
rect 512730 280412 512736 280424
rect 492088 280384 512736 280412
rect 492088 280372 492094 280384
rect 512730 280372 512736 280384
rect 512788 280372 512794 280424
rect 36998 280304 37004 280356
rect 37056 280344 37062 280356
rect 53650 280344 53656 280356
rect 37056 280316 53656 280344
rect 37056 280304 37062 280316
rect 53650 280304 53656 280316
rect 53708 280304 53714 280356
rect 148410 280304 148416 280356
rect 148468 280344 148474 280356
rect 165706 280344 165712 280356
rect 148468 280316 165712 280344
rect 148468 280304 148474 280316
rect 165706 280304 165712 280316
rect 165764 280304 165770 280356
rect 175458 280304 175464 280356
rect 175516 280344 175522 280356
rect 193674 280344 193680 280356
rect 175516 280316 193680 280344
rect 175516 280304 175522 280316
rect 193674 280304 193680 280316
rect 193732 280304 193738 280356
rect 203518 280304 203524 280356
rect 203576 280344 203582 280356
rect 221366 280344 221372 280356
rect 203576 280316 221372 280344
rect 203576 280304 203582 280316
rect 221366 280304 221372 280316
rect 221424 280304 221430 280356
rect 260098 280304 260104 280356
rect 260156 280344 260162 280356
rect 277670 280344 277676 280356
rect 260156 280316 277676 280344
rect 260156 280304 260162 280316
rect 277670 280304 277676 280316
rect 277728 280304 277734 280356
rect 287514 280304 287520 280356
rect 287572 280344 287578 280356
rect 305362 280344 305368 280356
rect 287572 280316 305368 280344
rect 287572 280304 287578 280316
rect 305362 280304 305368 280316
rect 305420 280304 305426 280356
rect 345658 280304 345664 280356
rect 345716 280344 345722 280356
rect 361666 280344 361672 280356
rect 345716 280316 361672 280344
rect 345716 280304 345722 280316
rect 361666 280304 361672 280316
rect 361724 280304 361730 280356
rect 371510 280304 371516 280356
rect 371568 280344 371574 280356
rect 389358 280344 389364 280356
rect 371568 280316 389364 280344
rect 371568 280304 371574 280316
rect 389358 280304 389364 280316
rect 389416 280304 389422 280356
rect 399478 280304 399484 280356
rect 399536 280344 399542 280356
rect 417694 280344 417700 280356
rect 399536 280316 417700 280344
rect 399536 280304 399542 280316
rect 417694 280304 417700 280316
rect 417752 280304 417758 280356
rect 456150 280304 456156 280356
rect 456208 280344 456214 280356
rect 473354 280344 473360 280356
rect 456208 280316 473360 280344
rect 456208 280304 456214 280316
rect 473354 280304 473360 280316
rect 473412 280304 473418 280356
rect 483474 280304 483480 280356
rect 483532 280344 483538 280356
rect 501690 280344 501696 280356
rect 483532 280316 501696 280344
rect 483532 280304 483538 280316
rect 501690 280304 501696 280316
rect 501748 280304 501754 280356
rect 36906 280236 36912 280288
rect 36964 280276 36970 280288
rect 63310 280276 63316 280288
rect 36964 280248 63316 280276
rect 36964 280236 36970 280248
rect 63310 280236 63316 280248
rect 63368 280236 63374 280288
rect 64322 280236 64328 280288
rect 64380 280276 64386 280288
rect 81434 280276 81440 280288
rect 64380 280248 81440 280276
rect 64380 280236 64386 280248
rect 81434 280236 81440 280248
rect 81492 280236 81498 280288
rect 91462 280236 91468 280288
rect 91520 280276 91526 280288
rect 109678 280276 109684 280288
rect 91520 280248 109684 280276
rect 91520 280236 91526 280248
rect 109678 280236 109684 280248
rect 109736 280236 109742 280288
rect 119430 280236 119436 280288
rect 119488 280276 119494 280288
rect 137646 280276 137652 280288
rect 119488 280248 137652 280276
rect 119488 280236 119494 280248
rect 137646 280236 137652 280248
rect 137704 280236 137710 280288
rect 156322 280236 156328 280288
rect 156380 280276 156386 280288
rect 178678 280276 178684 280288
rect 156380 280248 178684 280276
rect 156380 280236 156386 280248
rect 178678 280236 178684 280248
rect 178736 280236 178742 280288
rect 232498 280236 232504 280288
rect 232556 280276 232562 280288
rect 249702 280276 249708 280288
rect 232556 280248 249708 280276
rect 232556 280236 232562 280248
rect 249702 280236 249708 280248
rect 249760 280236 249766 280288
rect 268010 280236 268016 280288
rect 268068 280276 268074 280288
rect 287698 280276 287704 280288
rect 268068 280248 287704 280276
rect 268068 280236 268074 280248
rect 287698 280236 287704 280248
rect 287756 280236 287762 280288
rect 315482 280236 315488 280288
rect 315540 280276 315546 280288
rect 333698 280276 333704 280288
rect 315540 280248 333704 280276
rect 315540 280236 315546 280248
rect 333698 280236 333704 280248
rect 333756 280236 333762 280288
rect 352006 280236 352012 280288
rect 352064 280276 352070 280288
rect 374638 280276 374644 280288
rect 352064 280248 374644 280276
rect 352064 280236 352070 280248
rect 374638 280236 374644 280248
rect 374696 280236 374702 280288
rect 428458 280236 428464 280288
rect 428516 280276 428522 280288
rect 445662 280276 445668 280288
rect 428516 280248 445668 280276
rect 428516 280236 428522 280248
rect 445662 280236 445668 280248
rect 445720 280236 445726 280288
rect 464338 280236 464344 280288
rect 464396 280276 464402 280288
rect 483658 280276 483664 280288
rect 464396 280248 483664 280276
rect 464396 280236 464402 280248
rect 483658 280236 483664 280248
rect 483716 280236 483722 280288
rect 511442 280236 511448 280288
rect 511500 280276 511506 280288
rect 529658 280276 529664 280288
rect 511500 280248 529664 280276
rect 511500 280236 511506 280248
rect 529658 280236 529664 280248
rect 529716 280236 529722 280288
rect 542998 280236 543004 280288
rect 543056 280276 543062 280288
rect 557534 280276 557540 280288
rect 543056 280248 557540 280276
rect 543056 280236 543062 280248
rect 557534 280236 557540 280248
rect 557592 280236 557598 280288
rect 69658 280168 69664 280220
rect 69716 280208 69722 280220
rect 91094 280208 91100 280220
rect 69716 280180 91100 280208
rect 69716 280168 69722 280180
rect 91094 280168 91100 280180
rect 91152 280168 91158 280220
rect 94498 280168 94504 280220
rect 94556 280208 94562 280220
rect 119338 280208 119344 280220
rect 94556 280180 119344 280208
rect 94556 280168 94562 280180
rect 119338 280168 119344 280180
rect 119396 280168 119402 280220
rect 120718 280168 120724 280220
rect 120776 280208 120782 280220
rect 147306 280208 147312 280220
rect 120776 280180 147312 280208
rect 120776 280168 120782 280180
rect 147306 280168 147312 280180
rect 147364 280168 147370 280220
rect 148318 280168 148324 280220
rect 148376 280208 148382 280220
rect 175366 280208 175372 280220
rect 148376 280180 175372 280208
rect 148376 280168 148382 280180
rect 175366 280168 175372 280180
rect 175424 280168 175430 280220
rect 177298 280168 177304 280220
rect 177356 280208 177362 280220
rect 203334 280208 203340 280220
rect 177356 280180 203340 280208
rect 177356 280168 177362 280180
rect 203334 280168 203340 280180
rect 203392 280168 203398 280220
rect 204898 280168 204904 280220
rect 204956 280208 204962 280220
rect 231026 280208 231032 280220
rect 204956 280180 231032 280208
rect 204956 280168 204962 280180
rect 231026 280168 231032 280180
rect 231084 280168 231090 280220
rect 232590 280168 232596 280220
rect 232648 280208 232654 280220
rect 259362 280208 259368 280220
rect 232648 280180 259368 280208
rect 232648 280168 232654 280180
rect 259362 280168 259368 280180
rect 259420 280168 259426 280220
rect 260190 280168 260196 280220
rect 260248 280208 260254 280220
rect 287330 280208 287336 280220
rect 260248 280180 287336 280208
rect 260248 280168 260254 280180
rect 287330 280168 287336 280180
rect 287388 280168 287394 280220
rect 289078 280168 289084 280220
rect 289136 280208 289142 280220
rect 315022 280208 315028 280220
rect 289136 280180 315028 280208
rect 289136 280168 289142 280180
rect 315022 280168 315028 280180
rect 315080 280168 315086 280220
rect 316678 280168 316684 280220
rect 316736 280208 316742 280220
rect 343358 280208 343364 280220
rect 316736 280180 343364 280208
rect 316736 280168 316742 280180
rect 343358 280168 343364 280180
rect 343416 280168 343422 280220
rect 344278 280168 344284 280220
rect 344336 280208 344342 280220
rect 371326 280208 371332 280220
rect 344336 280180 371332 280208
rect 344336 280168 344342 280180
rect 371326 280168 371332 280180
rect 371384 280168 371390 280220
rect 373258 280168 373264 280220
rect 373316 280208 373322 280220
rect 399018 280208 399024 280220
rect 373316 280180 399024 280208
rect 373316 280168 373322 280180
rect 399018 280168 399024 280180
rect 399076 280168 399082 280220
rect 400858 280168 400864 280220
rect 400916 280208 400922 280220
rect 427354 280208 427360 280220
rect 400916 280180 427360 280208
rect 400916 280168 400922 280180
rect 427354 280168 427360 280180
rect 427412 280168 427418 280220
rect 428550 280168 428556 280220
rect 428608 280208 428614 280220
rect 455322 280208 455328 280220
rect 428608 280180 455328 280208
rect 428608 280168 428614 280180
rect 455322 280168 455328 280180
rect 455380 280168 455386 280220
rect 456058 280168 456064 280220
rect 456116 280208 456122 280220
rect 483014 280208 483020 280220
rect 456116 280180 483020 280208
rect 456116 280168 456122 280180
rect 483014 280168 483020 280180
rect 483072 280168 483078 280220
rect 485038 280168 485044 280220
rect 485096 280208 485102 280220
rect 511350 280208 511356 280220
rect 485096 280180 511356 280208
rect 485096 280168 485102 280180
rect 511350 280168 511356 280180
rect 511408 280168 511414 280220
rect 512638 280168 512644 280220
rect 512696 280208 512702 280220
rect 539318 280208 539324 280220
rect 512696 280180 539324 280208
rect 512696 280168 512702 280180
rect 539318 280168 539324 280180
rect 539376 280168 539382 280220
rect 540238 280168 540244 280220
rect 540296 280208 540302 280220
rect 567194 280208 567200 280220
rect 540296 280180 567200 280208
rect 540296 280168 540302 280180
rect 567194 280168 567200 280180
rect 567252 280168 567258 280220
rect 37918 279420 37924 279472
rect 37976 279460 37982 279472
rect 545758 279460 545764 279472
rect 37976 279432 545764 279460
rect 37976 279420 37982 279432
rect 545758 279420 545764 279432
rect 545816 279420 545822 279472
rect 182082 277516 182088 277568
rect 182140 277556 182146 277568
rect 233234 277556 233240 277568
rect 182140 277528 233240 277556
rect 182140 277516 182146 277528
rect 233234 277516 233240 277528
rect 233292 277516 233298 277568
rect 378042 277516 378048 277568
rect 378100 277556 378106 277568
rect 429194 277556 429200 277568
rect 378100 277528 429200 277556
rect 378100 277516 378106 277528
rect 429194 277516 429200 277528
rect 429252 277516 429258 277568
rect 462222 277516 462228 277568
rect 462280 277556 462286 277568
rect 513374 277556 513380 277568
rect 462280 277528 513380 277556
rect 462280 277516 462286 277528
rect 513374 277516 513380 277528
rect 513432 277516 513438 277568
rect 35618 277448 35624 277500
rect 35676 277488 35682 277500
rect 36814 277488 36820 277500
rect 35676 277460 36820 277488
rect 35676 277448 35682 277460
rect 36814 277448 36820 277460
rect 36872 277448 36878 277500
rect 42702 277448 42708 277500
rect 42760 277488 42766 277500
rect 93854 277488 93860 277500
rect 42760 277460 93860 277488
rect 42760 277448 42766 277460
rect 93854 277448 93860 277460
rect 93912 277448 93918 277500
rect 97902 277448 97908 277500
rect 97960 277488 97966 277500
rect 149054 277488 149060 277500
rect 97960 277460 149060 277488
rect 97960 277448 97966 277460
rect 149054 277448 149060 277460
rect 149112 277448 149118 277500
rect 154482 277448 154488 277500
rect 154540 277488 154546 277500
rect 205634 277488 205640 277500
rect 154540 277460 205640 277488
rect 154540 277448 154546 277460
rect 205634 277448 205640 277460
rect 205692 277448 205698 277500
rect 238662 277448 238668 277500
rect 238720 277488 238726 277500
rect 289814 277488 289820 277500
rect 238720 277460 289820 277488
rect 238720 277448 238726 277460
rect 289814 277448 289820 277460
rect 289872 277448 289878 277500
rect 293862 277448 293868 277500
rect 293920 277488 293926 277500
rect 345014 277488 345020 277500
rect 293920 277460 345020 277488
rect 293920 277448 293926 277460
rect 345014 277448 345020 277460
rect 345072 277448 345078 277500
rect 350442 277448 350448 277500
rect 350500 277488 350506 277500
rect 401594 277488 401600 277500
rect 350500 277460 401600 277488
rect 350500 277448 350506 277460
rect 401594 277448 401600 277460
rect 401652 277448 401658 277500
rect 434622 277448 434628 277500
rect 434680 277488 434686 277500
rect 485774 277488 485780 277500
rect 434680 277460 485780 277488
rect 434680 277448 434686 277460
rect 485774 277448 485780 277460
rect 485832 277448 485838 277500
rect 518802 277448 518808 277500
rect 518860 277488 518866 277500
rect 569954 277488 569960 277500
rect 518860 277460 569960 277488
rect 518860 277448 518866 277460
rect 569954 277448 569960 277460
rect 570012 277448 570018 277500
rect 13722 277380 13728 277432
rect 13780 277420 13786 277432
rect 66254 277420 66260 277432
rect 13780 277392 66260 277420
rect 13780 277380 13786 277392
rect 66254 277380 66260 277392
rect 66312 277380 66318 277432
rect 70302 277380 70308 277432
rect 70360 277420 70366 277432
rect 121454 277420 121460 277432
rect 70360 277392 121460 277420
rect 70360 277380 70366 277392
rect 121454 277380 121460 277392
rect 121512 277380 121518 277432
rect 126882 277380 126888 277432
rect 126940 277420 126946 277432
rect 178034 277420 178040 277432
rect 126940 277392 178040 277420
rect 126940 277380 126946 277392
rect 178034 277380 178040 277392
rect 178092 277380 178098 277432
rect 209682 277380 209688 277432
rect 209740 277420 209746 277432
rect 262214 277420 262220 277432
rect 209740 277392 262220 277420
rect 209740 277380 209746 277392
rect 262214 277380 262220 277392
rect 262272 277380 262278 277432
rect 266262 277380 266268 277432
rect 266320 277420 266326 277432
rect 317414 277420 317420 277432
rect 266320 277392 317420 277420
rect 266320 277380 266326 277392
rect 317414 277380 317420 277392
rect 317472 277380 317478 277432
rect 322842 277380 322848 277432
rect 322900 277420 322906 277432
rect 373994 277420 374000 277432
rect 322900 277392 374000 277420
rect 322900 277380 322906 277392
rect 373994 277380 374000 277392
rect 374052 277380 374058 277432
rect 405642 277380 405648 277432
rect 405700 277420 405706 277432
rect 458174 277420 458180 277432
rect 405700 277392 458180 277420
rect 405700 277380 405706 277392
rect 458174 277380 458180 277392
rect 458232 277380 458238 277432
rect 489822 277380 489828 277432
rect 489880 277420 489886 277432
rect 542354 277420 542360 277432
rect 489880 277392 542360 277420
rect 489880 277380 489886 277392
rect 542354 277380 542360 277392
rect 542412 277380 542418 277432
rect 63586 263440 63592 263492
rect 63644 263480 63650 263492
rect 64322 263480 64328 263492
rect 63644 263452 64328 263480
rect 63644 263440 63650 263452
rect 64322 263440 64328 263452
rect 64380 263440 64386 263492
rect 455690 263440 455696 263492
rect 455748 263480 455754 263492
rect 456150 263480 456156 263492
rect 455748 263452 456156 263480
rect 455748 263440 455754 263452
rect 456150 263440 456156 263452
rect 456208 263440 456214 263492
rect 232682 262148 232688 262200
rect 232740 262188 232746 262200
rect 239766 262188 239772 262200
rect 232740 262160 239772 262188
rect 232740 262148 232746 262160
rect 239766 262148 239772 262160
rect 239824 262148 239830 262200
rect 483658 262148 483664 262200
rect 483716 262188 483722 262200
rect 491662 262188 491668 262200
rect 483716 262160 491668 262188
rect 483716 262148 483722 262160
rect 491662 262148 491668 262160
rect 491720 262148 491726 262200
rect 512730 262148 512736 262200
rect 512788 262188 512794 262200
rect 519630 262188 519636 262200
rect 512788 262160 519636 262188
rect 512788 262148 512794 262160
rect 519630 262148 519636 262160
rect 519688 262148 519694 262200
rect 428642 261468 428648 261520
rect 428700 261508 428706 261520
rect 435726 261508 435732 261520
rect 428700 261480 435732 261508
rect 428700 261468 428706 261480
rect 435726 261468 435732 261480
rect 435784 261468 435790 261520
rect 316770 261400 316776 261452
rect 316828 261440 316834 261452
rect 323670 261440 323676 261452
rect 316828 261412 323676 261440
rect 316828 261400 316834 261412
rect 323670 261400 323676 261412
rect 323728 261400 323734 261452
rect 287698 261264 287704 261316
rect 287756 261304 287762 261316
rect 295702 261304 295708 261316
rect 287756 261276 295708 261304
rect 287756 261264 287762 261276
rect 295702 261264 295708 261276
rect 295760 261264 295766 261316
rect 147674 259428 147680 259480
rect 147732 259468 147738 259480
rect 148410 259468 148416 259480
rect 147732 259440 148416 259468
rect 147732 259428 147738 259440
rect 148410 259428 148416 259440
rect 148468 259428 148474 259480
rect 35618 259360 35624 259412
rect 35676 259400 35682 259412
rect 36998 259400 37004 259412
rect 35676 259372 37004 259400
rect 35676 259360 35682 259372
rect 36998 259360 37004 259372
rect 37056 259360 37062 259412
rect 343634 259360 343640 259412
rect 343692 259400 343698 259412
rect 345658 259400 345664 259412
rect 343692 259372 345664 259400
rect 343692 259360 343698 259372
rect 345658 259360 345664 259372
rect 345716 259360 345722 259412
rect 42886 256640 42892 256692
rect 42944 256680 42950 256692
rect 71958 256680 71964 256692
rect 42944 256652 45554 256680
rect 42944 256640 42950 256652
rect 15194 256572 15200 256624
rect 15252 256612 15258 256624
rect 43990 256612 43996 256624
rect 15252 256584 43996 256612
rect 15252 256572 15258 256584
rect 43990 256572 43996 256584
rect 44048 256572 44054 256624
rect 45526 256612 45554 256652
rect 64846 256652 71964 256680
rect 64846 256612 64874 256652
rect 71958 256640 71964 256652
rect 72016 256640 72022 256692
rect 99466 256640 99472 256692
rect 99524 256680 99530 256692
rect 99524 256652 103514 256680
rect 99524 256640 99530 256652
rect 45526 256584 64874 256612
rect 71866 256572 71872 256624
rect 71924 256612 71930 256624
rect 100018 256612 100024 256624
rect 71924 256584 100024 256612
rect 71924 256572 71930 256584
rect 100018 256572 100024 256584
rect 100076 256572 100082 256624
rect 103486 256612 103514 256652
rect 127066 256640 127072 256692
rect 127124 256680 127130 256692
rect 127124 256652 132494 256680
rect 127124 256640 127130 256652
rect 127986 256612 127992 256624
rect 103486 256584 127992 256612
rect 127986 256572 127992 256584
rect 128044 256572 128050 256624
rect 132466 256612 132494 256652
rect 183646 256640 183652 256692
rect 183704 256680 183710 256692
rect 183704 256652 190454 256680
rect 183704 256640 183710 256652
rect 155954 256612 155960 256624
rect 132466 256584 155960 256612
rect 155954 256572 155960 256584
rect 156012 256572 156018 256624
rect 165982 256572 165988 256624
rect 166040 256612 166046 256624
rect 177298 256612 177304 256624
rect 166040 256584 177304 256612
rect 166040 256572 166046 256584
rect 177298 256572 177304 256584
rect 177356 256572 177362 256624
rect 178678 256572 178684 256624
rect 178736 256612 178742 256624
rect 184014 256612 184020 256624
rect 178736 256584 184020 256612
rect 178736 256572 178742 256584
rect 184014 256572 184020 256584
rect 184072 256572 184078 256624
rect 190426 256612 190454 256652
rect 374638 256640 374644 256692
rect 374696 256680 374702 256692
rect 379698 256680 379704 256692
rect 374696 256652 379704 256680
rect 374696 256640 374702 256652
rect 379698 256640 379704 256652
rect 379756 256640 379762 256692
rect 539318 256640 539324 256692
rect 539376 256680 539382 256692
rect 542998 256680 543004 256692
rect 539376 256652 543004 256680
rect 539376 256640 539382 256652
rect 542998 256640 543004 256652
rect 543056 256640 543062 256692
rect 211706 256612 211712 256624
rect 190426 256584 211712 256612
rect 211706 256572 211712 256584
rect 211764 256572 211770 256624
rect 221918 256572 221924 256624
rect 221976 256612 221982 256624
rect 232590 256612 232596 256624
rect 221976 256584 232596 256612
rect 221976 256572 221982 256584
rect 232590 256572 232596 256584
rect 232648 256572 232654 256624
rect 249702 256572 249708 256624
rect 249760 256612 249766 256624
rect 260190 256612 260196 256624
rect 249760 256584 260196 256612
rect 249760 256572 249766 256584
rect 260190 256572 260196 256584
rect 260248 256572 260254 256624
rect 261478 256572 261484 256624
rect 261536 256612 261542 256624
rect 567194 256612 567200 256624
rect 261536 256584 567200 256612
rect 261536 256572 261542 256584
rect 567194 256572 567200 256584
rect 567252 256572 567258 256624
rect 25682 256504 25688 256556
rect 25740 256544 25746 256556
rect 36906 256544 36912 256556
rect 25740 256516 36912 256544
rect 25740 256504 25746 256516
rect 36906 256504 36912 256516
rect 36964 256504 36970 256556
rect 53650 256504 53656 256556
rect 53708 256544 53714 256556
rect 69658 256544 69664 256556
rect 53708 256516 69664 256544
rect 53708 256504 53714 256516
rect 69658 256504 69664 256516
rect 69716 256504 69722 256556
rect 81986 256504 81992 256556
rect 82044 256544 82050 256556
rect 94498 256544 94504 256556
rect 82044 256516 94504 256544
rect 82044 256504 82050 256516
rect 94498 256504 94504 256516
rect 94556 256504 94562 256556
rect 109678 256504 109684 256556
rect 109736 256544 109742 256556
rect 120718 256544 120724 256556
rect 109736 256516 120724 256544
rect 109736 256504 109742 256516
rect 120718 256504 120724 256516
rect 120776 256504 120782 256556
rect 137646 256504 137652 256556
rect 137704 256544 137710 256556
rect 148318 256544 148324 256556
rect 137704 256516 148324 256544
rect 137704 256504 137710 256516
rect 148318 256504 148324 256516
rect 148376 256504 148382 256556
rect 193674 256504 193680 256556
rect 193732 256544 193738 256556
rect 204898 256544 204904 256556
rect 193732 256516 204904 256544
rect 193732 256504 193738 256516
rect 204898 256504 204904 256516
rect 204956 256504 204962 256556
rect 238846 256504 238852 256556
rect 238904 256544 238910 256556
rect 268010 256544 268016 256556
rect 238904 256516 268016 256544
rect 238904 256504 238910 256516
rect 268010 256504 268016 256516
rect 268068 256504 268074 256556
rect 277670 256504 277676 256556
rect 277728 256544 277734 256556
rect 289078 256544 289084 256556
rect 277728 256516 289084 256544
rect 277728 256504 277734 256516
rect 289078 256504 289084 256516
rect 289136 256504 289142 256556
rect 306006 256504 306012 256556
rect 306064 256544 306070 256556
rect 316678 256544 316684 256556
rect 306064 256516 316684 256544
rect 306064 256504 306070 256516
rect 316678 256504 316684 256516
rect 316736 256504 316742 256556
rect 323026 256504 323032 256556
rect 323084 256544 323090 256556
rect 352006 256544 352012 256556
rect 323084 256516 352012 256544
rect 323084 256504 323090 256516
rect 352006 256504 352012 256516
rect 352064 256504 352070 256556
rect 361666 256504 361672 256556
rect 361724 256544 361730 256556
rect 373258 256544 373264 256556
rect 361724 256516 373264 256544
rect 361724 256504 361730 256516
rect 373258 256504 373264 256516
rect 373316 256504 373322 256556
rect 379606 256504 379612 256556
rect 379664 256544 379670 256556
rect 408034 256544 408040 256556
rect 379664 256516 408040 256544
rect 379664 256504 379670 256516
rect 408034 256504 408040 256516
rect 408092 256504 408098 256556
rect 417694 256504 417700 256556
rect 417752 256544 417758 256556
rect 428550 256544 428556 256556
rect 417752 256516 428556 256544
rect 417752 256504 417758 256516
rect 428550 256504 428556 256516
rect 428608 256504 428614 256556
rect 434806 256504 434812 256556
rect 434864 256544 434870 256556
rect 463786 256544 463792 256556
rect 434864 256516 463792 256544
rect 434864 256504 434870 256516
rect 463786 256504 463792 256516
rect 463844 256504 463850 256556
rect 473998 256504 474004 256556
rect 474056 256544 474062 256556
rect 485038 256544 485044 256556
rect 474056 256516 485044 256544
rect 474056 256504 474062 256516
rect 485038 256504 485044 256516
rect 485096 256504 485102 256556
rect 501690 256504 501696 256556
rect 501748 256544 501754 256556
rect 512638 256544 512644 256556
rect 501748 256516 512644 256544
rect 501748 256504 501754 256516
rect 512638 256504 512644 256516
rect 512696 256504 512702 256556
rect 518986 256504 518992 256556
rect 519044 256544 519050 256556
rect 547874 256544 547880 256556
rect 519044 256516 547880 256544
rect 519044 256504 519050 256516
rect 547874 256504 547880 256516
rect 547932 256504 547938 256556
rect 333698 256436 333704 256488
rect 333756 256476 333762 256488
rect 344278 256476 344284 256488
rect 333756 256448 344284 256476
rect 333756 256436 333762 256448
rect 344278 256436 344284 256448
rect 344336 256436 344342 256488
rect 390002 256436 390008 256488
rect 390060 256476 390066 256488
rect 400858 256476 400864 256488
rect 390060 256448 400864 256476
rect 390060 256436 390066 256448
rect 400858 256436 400864 256448
rect 400916 256436 400922 256488
rect 445662 256436 445668 256488
rect 445720 256476 445726 256488
rect 456058 256476 456064 256488
rect 445720 256448 456064 256476
rect 445720 256436 445726 256448
rect 456058 256436 456064 256448
rect 456116 256436 456122 256488
rect 529658 256436 529664 256488
rect 529716 256476 529722 256488
rect 540238 256476 540244 256488
rect 529716 256448 540244 256476
rect 529716 256436 529722 256448
rect 540238 256436 540244 256448
rect 540296 256436 540302 256488
rect 36722 256368 36728 256420
rect 36780 256408 36786 256420
rect 557534 256408 557540 256420
rect 36780 256380 557540 256408
rect 36780 256368 36786 256380
rect 557534 256368 557540 256380
rect 557592 256368 557598 256420
rect 16022 254532 16028 254584
rect 16080 254572 16086 254584
rect 547874 254572 547880 254584
rect 16080 254544 547880 254572
rect 16080 254532 16086 254544
rect 547874 254532 547880 254544
rect 547932 254532 547938 254584
rect 25682 254124 25688 254176
rect 25740 254164 25746 254176
rect 69658 254164 69664 254176
rect 25740 254136 69664 254164
rect 25740 254124 25746 254136
rect 69658 254124 69664 254136
rect 69716 254124 69722 254176
rect 212350 254124 212356 254176
rect 212408 254164 212414 254176
rect 232682 254164 232688 254176
rect 212408 254136 232688 254164
rect 212408 254124 212414 254136
rect 232682 254124 232688 254136
rect 232740 254124 232746 254176
rect 296346 254124 296352 254176
rect 296404 254164 296410 254176
rect 316770 254164 316776 254176
rect 296404 254136 316776 254164
rect 296404 254124 296410 254136
rect 316770 254124 316776 254136
rect 316828 254124 316834 254176
rect 492030 254124 492036 254176
rect 492088 254164 492094 254176
rect 512730 254164 512736 254176
rect 492088 254136 512736 254164
rect 492088 254124 492094 254136
rect 512730 254124 512736 254136
rect 512788 254124 512794 254176
rect 3326 254056 3332 254108
rect 3384 254096 3390 254108
rect 7650 254096 7656 254108
rect 3384 254068 7656 254096
rect 3384 254056 3390 254068
rect 7650 254056 7656 254068
rect 7708 254056 7714 254108
rect 36998 254056 37004 254108
rect 37056 254096 37062 254108
rect 53650 254096 53656 254108
rect 37056 254068 53656 254096
rect 37056 254056 37062 254068
rect 53650 254056 53656 254068
rect 53708 254056 53714 254108
rect 64322 254056 64328 254108
rect 64380 254096 64386 254108
rect 81434 254096 81440 254108
rect 64380 254068 81440 254096
rect 64380 254056 64386 254068
rect 81434 254056 81440 254068
rect 81492 254056 81498 254108
rect 148410 254056 148416 254108
rect 148468 254096 148474 254108
rect 165706 254096 165712 254108
rect 148468 254068 165712 254096
rect 148468 254056 148474 254068
rect 165706 254056 165712 254068
rect 165764 254056 165770 254108
rect 175458 254056 175464 254108
rect 175516 254096 175522 254108
rect 193674 254096 193680 254108
rect 175516 254068 193680 254096
rect 175516 254056 175522 254068
rect 193674 254056 193680 254068
rect 193732 254056 193738 254108
rect 203518 254056 203524 254108
rect 203576 254096 203582 254108
rect 221366 254096 221372 254108
rect 203576 254068 221372 254096
rect 203576 254056 203582 254068
rect 221366 254056 221372 254068
rect 221424 254056 221430 254108
rect 260190 254056 260196 254108
rect 260248 254096 260254 254108
rect 277670 254096 277676 254108
rect 260248 254068 277676 254096
rect 260248 254056 260254 254068
rect 277670 254056 277676 254068
rect 277728 254056 277734 254108
rect 287514 254056 287520 254108
rect 287572 254096 287578 254108
rect 305362 254096 305368 254108
rect 287572 254068 305368 254096
rect 287572 254056 287578 254068
rect 305362 254056 305368 254068
rect 305420 254056 305426 254108
rect 345658 254056 345664 254108
rect 345716 254096 345722 254108
rect 361666 254096 361672 254108
rect 345716 254068 361672 254096
rect 345716 254056 345722 254068
rect 361666 254056 361672 254068
rect 361724 254056 361730 254108
rect 371510 254056 371516 254108
rect 371568 254096 371574 254108
rect 389358 254096 389364 254108
rect 371568 254068 389364 254096
rect 371568 254056 371574 254068
rect 389358 254056 389364 254068
rect 389416 254056 389422 254108
rect 399478 254056 399484 254108
rect 399536 254096 399542 254108
rect 417694 254096 417700 254108
rect 399536 254068 417700 254096
rect 399536 254056 399542 254068
rect 417694 254056 417700 254068
rect 417752 254056 417758 254108
rect 428550 254056 428556 254108
rect 428608 254096 428614 254108
rect 445662 254096 445668 254108
rect 428608 254068 445668 254096
rect 428608 254056 428614 254068
rect 445662 254056 445668 254068
rect 445720 254056 445726 254108
rect 456058 254056 456064 254108
rect 456116 254096 456122 254108
rect 473354 254096 473360 254108
rect 456116 254068 473360 254096
rect 456116 254056 456122 254068
rect 473354 254056 473360 254068
rect 473412 254056 473418 254108
rect 483474 254056 483480 254108
rect 483532 254096 483538 254108
rect 501690 254096 501696 254108
rect 483532 254068 501696 254096
rect 483532 254056 483538 254068
rect 501690 254056 501696 254068
rect 501748 254056 501754 254108
rect 36906 253988 36912 254040
rect 36964 254028 36970 254040
rect 63310 254028 63316 254040
rect 36964 254000 63316 254028
rect 36964 253988 36970 254000
rect 63310 253988 63316 254000
rect 63368 253988 63374 254040
rect 66898 253988 66904 254040
rect 66956 254028 66962 254040
rect 91094 254028 91100 254040
rect 66956 254000 91100 254028
rect 66956 253988 66962 254000
rect 91094 253988 91100 254000
rect 91152 253988 91158 254040
rect 91462 253988 91468 254040
rect 91520 254028 91526 254040
rect 109678 254028 109684 254040
rect 91520 254000 109684 254028
rect 91520 253988 91526 254000
rect 109678 253988 109684 254000
rect 109736 253988 109742 254040
rect 119430 253988 119436 254040
rect 119488 254028 119494 254040
rect 137646 254028 137652 254040
rect 119488 254000 137652 254028
rect 119488 253988 119494 254000
rect 137646 253988 137652 254000
rect 137704 253988 137710 254040
rect 156322 253988 156328 254040
rect 156380 254028 156386 254040
rect 178678 254028 178684 254040
rect 156380 254000 178684 254028
rect 156380 253988 156386 254000
rect 178678 253988 178684 254000
rect 178736 253988 178742 254040
rect 232590 253988 232596 254040
rect 232648 254028 232654 254040
rect 249702 254028 249708 254040
rect 232648 254000 249708 254028
rect 232648 253988 232654 254000
rect 249702 253988 249708 254000
rect 249760 253988 249766 254040
rect 268010 253988 268016 254040
rect 268068 254028 268074 254040
rect 287698 254028 287704 254040
rect 268068 254000 287704 254028
rect 268068 253988 268074 254000
rect 287698 253988 287704 254000
rect 287756 253988 287762 254040
rect 315482 253988 315488 254040
rect 315540 254028 315546 254040
rect 333698 254028 333704 254040
rect 315540 254000 333704 254028
rect 315540 253988 315546 254000
rect 333698 253988 333704 254000
rect 333756 253988 333762 254040
rect 352006 253988 352012 254040
rect 352064 254028 352070 254040
rect 374638 254028 374644 254040
rect 352064 254000 374644 254028
rect 352064 253988 352070 254000
rect 374638 253988 374644 254000
rect 374696 253988 374702 254040
rect 408034 253988 408040 254040
rect 408092 254028 408098 254040
rect 428642 254028 428648 254040
rect 408092 254000 428648 254028
rect 408092 253988 408098 254000
rect 428642 253988 428648 254000
rect 428700 253988 428706 254040
rect 464338 253988 464344 254040
rect 464396 254028 464402 254040
rect 483658 254028 483664 254040
rect 464396 254000 483664 254028
rect 464396 253988 464402 254000
rect 483658 253988 483664 254000
rect 483716 253988 483722 254040
rect 511442 253988 511448 254040
rect 511500 254028 511506 254040
rect 529658 254028 529664 254040
rect 511500 254000 529664 254028
rect 511500 253988 511506 254000
rect 529658 253988 529664 254000
rect 529716 253988 529722 254040
rect 542998 253988 543004 254040
rect 543056 254028 543062 254040
rect 557534 254028 557540 254040
rect 543056 254000 557540 254028
rect 543056 253988 543062 254000
rect 557534 253988 557540 254000
rect 557592 253988 557598 254040
rect 94498 253920 94504 253972
rect 94556 253960 94562 253972
rect 119338 253960 119344 253972
rect 94556 253932 119344 253960
rect 94556 253920 94562 253932
rect 119338 253920 119344 253932
rect 119396 253920 119402 253972
rect 120718 253920 120724 253972
rect 120776 253960 120782 253972
rect 147306 253960 147312 253972
rect 120776 253932 147312 253960
rect 120776 253920 120782 253932
rect 147306 253920 147312 253932
rect 147364 253920 147370 253972
rect 148318 253920 148324 253972
rect 148376 253960 148382 253972
rect 175366 253960 175372 253972
rect 148376 253932 175372 253960
rect 148376 253920 148382 253932
rect 175366 253920 175372 253932
rect 175424 253920 175430 253972
rect 177298 253920 177304 253972
rect 177356 253960 177362 253972
rect 203334 253960 203340 253972
rect 177356 253932 203340 253960
rect 177356 253920 177362 253932
rect 203334 253920 203340 253932
rect 203392 253920 203398 253972
rect 204898 253920 204904 253972
rect 204956 253960 204962 253972
rect 231026 253960 231032 253972
rect 204956 253932 231032 253960
rect 204956 253920 204962 253932
rect 231026 253920 231032 253932
rect 231084 253920 231090 253972
rect 232498 253920 232504 253972
rect 232556 253960 232562 253972
rect 259362 253960 259368 253972
rect 232556 253932 259368 253960
rect 232556 253920 232562 253932
rect 259362 253920 259368 253932
rect 259420 253920 259426 253972
rect 260098 253920 260104 253972
rect 260156 253960 260162 253972
rect 287330 253960 287336 253972
rect 260156 253932 287336 253960
rect 260156 253920 260162 253932
rect 287330 253920 287336 253932
rect 287388 253920 287394 253972
rect 289078 253920 289084 253972
rect 289136 253960 289142 253972
rect 315022 253960 315028 253972
rect 289136 253932 315028 253960
rect 289136 253920 289142 253932
rect 315022 253920 315028 253932
rect 315080 253920 315086 253972
rect 316678 253920 316684 253972
rect 316736 253960 316742 253972
rect 343358 253960 343364 253972
rect 316736 253932 343364 253960
rect 316736 253920 316742 253932
rect 343358 253920 343364 253932
rect 343416 253920 343422 253972
rect 344278 253920 344284 253972
rect 344336 253960 344342 253972
rect 371326 253960 371332 253972
rect 344336 253932 371332 253960
rect 344336 253920 344342 253932
rect 371326 253920 371332 253932
rect 371384 253920 371390 253972
rect 373258 253920 373264 253972
rect 373316 253960 373322 253972
rect 399018 253960 399024 253972
rect 373316 253932 399024 253960
rect 373316 253920 373322 253932
rect 399018 253920 399024 253932
rect 399076 253920 399082 253972
rect 400858 253920 400864 253972
rect 400916 253960 400922 253972
rect 427354 253960 427360 253972
rect 400916 253932 427360 253960
rect 400916 253920 400922 253932
rect 427354 253920 427360 253932
rect 427412 253920 427418 253972
rect 428458 253920 428464 253972
rect 428516 253960 428522 253972
rect 455322 253960 455328 253972
rect 428516 253932 455328 253960
rect 428516 253920 428522 253932
rect 455322 253920 455328 253932
rect 455380 253920 455386 253972
rect 456150 253920 456156 253972
rect 456208 253960 456214 253972
rect 483014 253960 483020 253972
rect 456208 253932 483020 253960
rect 456208 253920 456214 253932
rect 483014 253920 483020 253932
rect 483072 253920 483078 253972
rect 485038 253920 485044 253972
rect 485096 253960 485102 253972
rect 511350 253960 511356 253972
rect 485096 253932 511356 253960
rect 485096 253920 485102 253932
rect 511350 253920 511356 253932
rect 511408 253920 511414 253972
rect 512638 253920 512644 253972
rect 512696 253960 512702 253972
rect 539318 253960 539324 253972
rect 512696 253932 539324 253960
rect 512696 253920 512702 253932
rect 539318 253920 539324 253932
rect 539376 253920 539382 253972
rect 540238 253920 540244 253972
rect 540296 253960 540302 253972
rect 567194 253960 567200 253972
rect 540296 253932 567200 253960
rect 540296 253920 540302 253932
rect 567194 253920 567200 253932
rect 567252 253920 567258 253972
rect 37918 251812 37924 251864
rect 37976 251852 37982 251864
rect 545758 251852 545764 251864
rect 37976 251824 545764 251852
rect 37976 251812 37982 251824
rect 545758 251812 545764 251824
rect 545816 251812 545822 251864
rect 182082 251268 182088 251320
rect 182140 251308 182146 251320
rect 233234 251308 233240 251320
rect 182140 251280 233240 251308
rect 182140 251268 182146 251280
rect 233234 251268 233240 251280
rect 233292 251268 233298 251320
rect 378042 251268 378048 251320
rect 378100 251308 378106 251320
rect 429194 251308 429200 251320
rect 378100 251280 429200 251308
rect 378100 251268 378106 251280
rect 429194 251268 429200 251280
rect 429252 251268 429258 251320
rect 35618 251200 35624 251252
rect 35676 251240 35682 251252
rect 36722 251240 36728 251252
rect 35676 251212 36728 251240
rect 35676 251200 35682 251212
rect 36722 251200 36728 251212
rect 36780 251200 36786 251252
rect 42702 251200 42708 251252
rect 42760 251240 42766 251252
rect 93854 251240 93860 251252
rect 42760 251212 93860 251240
rect 42760 251200 42766 251212
rect 93854 251200 93860 251212
rect 93912 251200 93918 251252
rect 97902 251200 97908 251252
rect 97960 251240 97966 251252
rect 149054 251240 149060 251252
rect 97960 251212 149060 251240
rect 97960 251200 97966 251212
rect 149054 251200 149060 251212
rect 149112 251200 149118 251252
rect 154482 251200 154488 251252
rect 154540 251240 154546 251252
rect 205634 251240 205640 251252
rect 154540 251212 205640 251240
rect 154540 251200 154546 251212
rect 205634 251200 205640 251212
rect 205692 251200 205698 251252
rect 238662 251200 238668 251252
rect 238720 251240 238726 251252
rect 289814 251240 289820 251252
rect 238720 251212 289820 251240
rect 238720 251200 238726 251212
rect 289814 251200 289820 251212
rect 289872 251200 289878 251252
rect 293862 251200 293868 251252
rect 293920 251240 293926 251252
rect 345014 251240 345020 251252
rect 293920 251212 345020 251240
rect 293920 251200 293926 251212
rect 345014 251200 345020 251212
rect 345072 251200 345078 251252
rect 350442 251200 350448 251252
rect 350500 251240 350506 251252
rect 401594 251240 401600 251252
rect 350500 251212 401600 251240
rect 350500 251200 350506 251212
rect 401594 251200 401600 251212
rect 401652 251200 401658 251252
rect 434622 251200 434628 251252
rect 434680 251240 434686 251252
rect 485774 251240 485780 251252
rect 434680 251212 485780 251240
rect 434680 251200 434686 251212
rect 485774 251200 485780 251212
rect 485832 251200 485838 251252
rect 489822 251200 489828 251252
rect 489880 251240 489886 251252
rect 542354 251240 542360 251252
rect 489880 251212 542360 251240
rect 489880 251200 489886 251212
rect 542354 251200 542360 251212
rect 542412 251200 542418 251252
rect 3050 240184 3056 240236
rect 3108 240224 3114 240236
rect 6270 240224 6276 240236
rect 3108 240196 6276 240224
rect 3108 240184 3114 240196
rect 6270 240184 6276 240196
rect 6328 240184 6334 240236
rect 63586 235356 63592 235408
rect 63644 235396 63650 235408
rect 64322 235396 64328 235408
rect 63644 235368 64328 235396
rect 63644 235356 63650 235368
rect 64322 235356 64328 235368
rect 64380 235356 64386 235408
rect 147674 235356 147680 235408
rect 147732 235396 147738 235408
rect 148410 235396 148416 235408
rect 147732 235368 148416 235396
rect 147732 235356 147738 235368
rect 148410 235356 148416 235368
rect 148468 235356 148474 235408
rect 259730 235356 259736 235408
rect 259788 235396 259794 235408
rect 260190 235396 260196 235408
rect 259788 235368 260196 235396
rect 259788 235356 259794 235368
rect 260190 235356 260196 235368
rect 260248 235356 260254 235408
rect 512730 234200 512736 234252
rect 512788 234240 512794 234252
rect 519630 234240 519636 234252
rect 512788 234212 519636 234240
rect 512788 234200 512794 234212
rect 519630 234200 519636 234212
rect 519688 234200 519694 234252
rect 428642 233860 428648 233912
rect 428700 233900 428706 233912
rect 435726 233900 435732 233912
rect 428700 233872 435732 233900
rect 428700 233860 428706 233872
rect 435726 233860 435732 233872
rect 435784 233860 435790 233912
rect 232682 233520 232688 233572
rect 232740 233560 232746 233572
rect 239766 233560 239772 233572
rect 232740 233532 239772 233560
rect 232740 233520 232746 233532
rect 239766 233520 239772 233532
rect 239824 233520 239830 233572
rect 287698 233520 287704 233572
rect 287756 233560 287762 233572
rect 295702 233560 295708 233572
rect 287756 233532 295708 233560
rect 287756 233520 287762 233532
rect 295702 233520 295708 233532
rect 295760 233520 295766 233572
rect 316770 233384 316776 233436
rect 316828 233424 316834 233436
rect 323670 233424 323676 233436
rect 316828 233396 323676 233424
rect 316828 233384 316834 233396
rect 323670 233384 323676 233396
rect 323728 233384 323734 233436
rect 483658 233384 483664 233436
rect 483716 233424 483722 233436
rect 491662 233424 491668 233436
rect 483716 233396 491668 233424
rect 483716 233384 483722 233396
rect 491662 233384 491668 233396
rect 491720 233384 491726 233436
rect 13722 233180 13728 233232
rect 13780 233220 13786 233232
rect 66254 233220 66260 233232
rect 13780 233192 66260 233220
rect 13780 233180 13786 233192
rect 66254 233180 66260 233192
rect 66312 233180 66318 233232
rect 70302 233180 70308 233232
rect 70360 233220 70366 233232
rect 121454 233220 121460 233232
rect 70360 233192 121460 233220
rect 70360 233180 70366 233192
rect 121454 233180 121460 233192
rect 121512 233180 121518 233232
rect 126882 233180 126888 233232
rect 126940 233220 126946 233232
rect 178034 233220 178040 233232
rect 126940 233192 178040 233220
rect 126940 233180 126946 233192
rect 178034 233180 178040 233192
rect 178092 233180 178098 233232
rect 209682 233180 209688 233232
rect 209740 233220 209746 233232
rect 262214 233220 262220 233232
rect 209740 233192 262220 233220
rect 209740 233180 209746 233192
rect 262214 233180 262220 233192
rect 262272 233180 262278 233232
rect 266262 233180 266268 233232
rect 266320 233220 266326 233232
rect 317414 233220 317420 233232
rect 266320 233192 317420 233220
rect 266320 233180 266326 233192
rect 317414 233180 317420 233192
rect 317472 233180 317478 233232
rect 322842 233180 322848 233232
rect 322900 233220 322906 233232
rect 373994 233220 374000 233232
rect 322900 233192 374000 233220
rect 322900 233180 322906 233192
rect 373994 233180 374000 233192
rect 374052 233180 374058 233232
rect 405642 233180 405648 233232
rect 405700 233220 405706 233232
rect 458174 233220 458180 233232
rect 405700 233192 458180 233220
rect 405700 233180 405706 233192
rect 458174 233180 458180 233192
rect 458232 233180 458238 233232
rect 462222 233180 462228 233232
rect 462280 233220 462286 233232
rect 513374 233220 513380 233232
rect 462280 233192 513380 233220
rect 462280 233180 462286 233192
rect 513374 233180 513380 233192
rect 513432 233180 513438 233232
rect 518802 233180 518808 233232
rect 518860 233220 518866 233232
rect 569954 233220 569960 233232
rect 518860 233192 569960 233220
rect 518860 233180 518866 233192
rect 569954 233180 569960 233192
rect 570012 233180 570018 233232
rect 231670 233112 231676 233164
rect 231728 233152 231734 233164
rect 232590 233152 232596 233164
rect 231728 233124 232596 233152
rect 231728 233112 231734 233124
rect 232590 233112 232596 233124
rect 232648 233112 232654 233164
rect 427722 233112 427728 233164
rect 427780 233152 427786 233164
rect 428550 233152 428556 233164
rect 427780 233124 428556 233152
rect 427780 233112 427786 233124
rect 428550 233112 428556 233124
rect 428608 233112 428614 233164
rect 539502 233112 539508 233164
rect 539560 233152 539566 233164
rect 542998 233152 543004 233164
rect 539560 233124 543004 233152
rect 539560 233112 539566 233124
rect 542998 233112 543004 233124
rect 543056 233112 543062 233164
rect 35618 232704 35624 232756
rect 35676 232744 35682 232756
rect 36998 232744 37004 232756
rect 35676 232716 37004 232744
rect 35676 232704 35682 232716
rect 36998 232704 37004 232716
rect 37056 232704 37062 232756
rect 343634 232704 343640 232756
rect 343692 232744 343698 232756
rect 345658 232744 345664 232756
rect 343692 232716 345664 232744
rect 343692 232704 343698 232716
rect 345658 232704 345664 232716
rect 345716 232704 345722 232756
rect 178678 230392 178684 230444
rect 178736 230432 178742 230444
rect 184014 230432 184020 230444
rect 178736 230404 184020 230432
rect 178736 230392 178742 230404
rect 184014 230392 184020 230404
rect 184072 230392 184078 230444
rect 374638 230392 374644 230444
rect 374696 230432 374702 230444
rect 379698 230432 379704 230444
rect 374696 230404 379704 230432
rect 374696 230392 374702 230404
rect 379698 230392 379704 230404
rect 379756 230392 379762 230444
rect 15194 230324 15200 230376
rect 15252 230364 15258 230376
rect 43990 230364 43996 230376
rect 15252 230336 43996 230364
rect 15252 230324 15258 230336
rect 43990 230324 43996 230336
rect 44048 230324 44054 230376
rect 71038 230324 71044 230376
rect 71096 230364 71102 230376
rect 567194 230364 567200 230376
rect 71096 230336 567200 230364
rect 71096 230324 71102 230336
rect 567194 230324 567200 230336
rect 567252 230324 567258 230376
rect 25682 230256 25688 230308
rect 25740 230296 25746 230308
rect 36906 230296 36912 230308
rect 25740 230268 36912 230296
rect 25740 230256 25746 230268
rect 36906 230256 36912 230268
rect 36964 230256 36970 230308
rect 53650 230256 53656 230308
rect 53708 230296 53714 230308
rect 66898 230296 66904 230308
rect 53708 230268 66904 230296
rect 53708 230256 53714 230268
rect 66898 230256 66904 230268
rect 66956 230256 66962 230308
rect 71866 230256 71872 230308
rect 71924 230296 71930 230308
rect 100018 230296 100024 230308
rect 71924 230268 100024 230296
rect 71924 230256 71930 230268
rect 100018 230256 100024 230268
rect 100076 230256 100082 230308
rect 127986 230296 127992 230308
rect 103486 230268 127992 230296
rect 42886 230188 42892 230240
rect 42944 230228 42950 230240
rect 72050 230228 72056 230240
rect 42944 230200 72056 230228
rect 42944 230188 42950 230200
rect 72050 230188 72056 230200
rect 72108 230188 72114 230240
rect 81986 230188 81992 230240
rect 82044 230228 82050 230240
rect 94498 230228 94504 230240
rect 82044 230200 94504 230228
rect 82044 230188 82050 230200
rect 94498 230188 94504 230200
rect 94556 230188 94562 230240
rect 99466 230188 99472 230240
rect 99524 230228 99530 230240
rect 103486 230228 103514 230268
rect 127986 230256 127992 230268
rect 128044 230256 128050 230308
rect 156046 230296 156052 230308
rect 132466 230268 156052 230296
rect 99524 230200 103514 230228
rect 99524 230188 99530 230200
rect 109678 230188 109684 230240
rect 109736 230228 109742 230240
rect 120718 230228 120724 230240
rect 109736 230200 120724 230228
rect 109736 230188 109742 230200
rect 120718 230188 120724 230200
rect 120776 230188 120782 230240
rect 127066 230188 127072 230240
rect 127124 230228 127130 230240
rect 132466 230228 132494 230268
rect 156046 230256 156052 230268
rect 156104 230256 156110 230308
rect 165982 230256 165988 230308
rect 166040 230296 166046 230308
rect 177298 230296 177304 230308
rect 166040 230268 177304 230296
rect 166040 230256 166046 230268
rect 177298 230256 177304 230268
rect 177356 230256 177362 230308
rect 183646 230256 183652 230308
rect 183704 230296 183710 230308
rect 211706 230296 211712 230308
rect 183704 230268 211712 230296
rect 183704 230256 183710 230268
rect 211706 230256 211712 230268
rect 211764 230256 211770 230308
rect 222010 230256 222016 230308
rect 222068 230296 222074 230308
rect 232498 230296 232504 230308
rect 222068 230268 232504 230296
rect 222068 230256 222074 230268
rect 232498 230256 232504 230268
rect 232556 230256 232562 230308
rect 238846 230256 238852 230308
rect 238904 230296 238910 230308
rect 268010 230296 268016 230308
rect 238904 230268 268016 230296
rect 238904 230256 238910 230268
rect 268010 230256 268016 230268
rect 268068 230256 268074 230308
rect 277670 230256 277676 230308
rect 277728 230296 277734 230308
rect 289078 230296 289084 230308
rect 277728 230268 289084 230296
rect 277728 230256 277734 230268
rect 289078 230256 289084 230268
rect 289136 230256 289142 230308
rect 306006 230256 306012 230308
rect 306064 230296 306070 230308
rect 316678 230296 316684 230308
rect 306064 230268 316684 230296
rect 306064 230256 306070 230268
rect 316678 230256 316684 230268
rect 316736 230256 316742 230308
rect 323026 230256 323032 230308
rect 323084 230296 323090 230308
rect 352006 230296 352012 230308
rect 323084 230268 352012 230296
rect 323084 230256 323090 230268
rect 352006 230256 352012 230268
rect 352064 230256 352070 230308
rect 361666 230256 361672 230308
rect 361724 230296 361730 230308
rect 373258 230296 373264 230308
rect 361724 230268 373264 230296
rect 361724 230256 361730 230268
rect 373258 230256 373264 230268
rect 373316 230256 373322 230308
rect 379606 230256 379612 230308
rect 379664 230296 379670 230308
rect 408034 230296 408040 230308
rect 379664 230268 408040 230296
rect 379664 230256 379670 230268
rect 408034 230256 408040 230268
rect 408092 230256 408098 230308
rect 417694 230256 417700 230308
rect 417752 230296 417758 230308
rect 428458 230296 428464 230308
rect 417752 230268 428464 230296
rect 417752 230256 417758 230268
rect 428458 230256 428464 230268
rect 428516 230256 428522 230308
rect 434806 230256 434812 230308
rect 434864 230296 434870 230308
rect 463694 230296 463700 230308
rect 434864 230268 463700 230296
rect 434864 230256 434870 230268
rect 463694 230256 463700 230268
rect 463752 230256 463758 230308
rect 473998 230256 474004 230308
rect 474056 230296 474062 230308
rect 485038 230296 485044 230308
rect 474056 230268 485044 230296
rect 474056 230256 474062 230268
rect 485038 230256 485044 230268
rect 485096 230256 485102 230308
rect 501690 230256 501696 230308
rect 501748 230296 501754 230308
rect 512638 230296 512644 230308
rect 501748 230268 512644 230296
rect 501748 230256 501754 230268
rect 512638 230256 512644 230268
rect 512696 230256 512702 230308
rect 518986 230256 518992 230308
rect 519044 230296 519050 230308
rect 547874 230296 547880 230308
rect 519044 230268 547880 230296
rect 519044 230256 519050 230268
rect 547874 230256 547880 230268
rect 547932 230256 547938 230308
rect 127124 230200 132494 230228
rect 127124 230188 127130 230200
rect 137646 230188 137652 230240
rect 137704 230228 137710 230240
rect 148318 230228 148324 230240
rect 137704 230200 148324 230228
rect 137704 230188 137710 230200
rect 148318 230188 148324 230200
rect 148376 230188 148382 230240
rect 193674 230188 193680 230240
rect 193732 230228 193738 230240
rect 204898 230228 204904 230240
rect 193732 230200 204904 230228
rect 193732 230188 193738 230200
rect 204898 230188 204904 230200
rect 204956 230188 204962 230240
rect 249702 230188 249708 230240
rect 249760 230228 249766 230240
rect 260098 230228 260104 230240
rect 249760 230200 260104 230228
rect 249760 230188 249766 230200
rect 260098 230188 260104 230200
rect 260156 230188 260162 230240
rect 333698 230188 333704 230240
rect 333756 230228 333762 230240
rect 344278 230228 344284 230240
rect 333756 230200 344284 230228
rect 333756 230188 333762 230200
rect 344278 230188 344284 230200
rect 344336 230188 344342 230240
rect 390002 230188 390008 230240
rect 390060 230228 390066 230240
rect 400858 230228 400864 230240
rect 390060 230200 400864 230228
rect 390060 230188 390066 230200
rect 400858 230188 400864 230200
rect 400916 230188 400922 230240
rect 445662 230188 445668 230240
rect 445720 230228 445726 230240
rect 456150 230228 456156 230240
rect 445720 230200 456156 230228
rect 445720 230188 445726 230200
rect 456150 230188 456156 230200
rect 456208 230188 456214 230240
rect 529658 230188 529664 230240
rect 529716 230228 529722 230240
rect 540238 230228 540244 230240
rect 529716 230200 540244 230228
rect 529716 230188 529722 230200
rect 540238 230188 540244 230200
rect 540296 230188 540302 230240
rect 36814 230120 36820 230172
rect 36872 230160 36878 230172
rect 557534 230160 557540 230172
rect 36872 230132 557540 230160
rect 36872 230120 36878 230132
rect 557534 230120 557540 230132
rect 557592 230120 557598 230172
rect 15286 226992 15292 227044
rect 15344 227032 15350 227044
rect 547874 227032 547880 227044
rect 15344 227004 547880 227032
rect 15344 226992 15350 227004
rect 547874 226992 547880 227004
rect 547932 226992 547938 227044
rect 25682 226584 25688 226636
rect 25740 226624 25746 226636
rect 261478 226624 261484 226636
rect 25740 226596 261484 226624
rect 25740 226584 25746 226596
rect 261478 226584 261484 226596
rect 261536 226584 261542 226636
rect 148318 226516 148324 226568
rect 148376 226556 148382 226568
rect 165706 226556 165712 226568
rect 148376 226528 165712 226556
rect 148376 226516 148382 226528
rect 165706 226516 165712 226528
rect 165764 226516 165770 226568
rect 175458 226516 175464 226568
rect 175516 226556 175522 226568
rect 193674 226556 193680 226568
rect 175516 226528 193680 226556
rect 175516 226516 175522 226528
rect 193674 226516 193680 226528
rect 193732 226516 193738 226568
rect 203518 226516 203524 226568
rect 203576 226556 203582 226568
rect 221366 226556 221372 226568
rect 203576 226528 221372 226556
rect 203576 226516 203582 226528
rect 221366 226516 221372 226528
rect 221424 226516 221430 226568
rect 296346 226516 296352 226568
rect 296404 226556 296410 226568
rect 316770 226556 316776 226568
rect 296404 226528 316776 226556
rect 296404 226516 296410 226528
rect 316770 226516 316776 226528
rect 316828 226516 316834 226568
rect 408034 226516 408040 226568
rect 408092 226556 408098 226568
rect 428642 226556 428648 226568
rect 408092 226528 428648 226556
rect 408092 226516 408098 226528
rect 428642 226516 428648 226528
rect 428700 226516 428706 226568
rect 492030 226516 492036 226568
rect 492088 226556 492094 226568
rect 512730 226556 512736 226568
rect 492088 226528 512736 226556
rect 492088 226516 492094 226528
rect 512730 226516 512736 226528
rect 512788 226516 512794 226568
rect 36998 226448 37004 226500
rect 37056 226488 37062 226500
rect 53650 226488 53656 226500
rect 37056 226460 53656 226488
rect 37056 226448 37062 226460
rect 53650 226448 53656 226460
rect 53708 226448 53714 226500
rect 64322 226448 64328 226500
rect 64380 226488 64386 226500
rect 81434 226488 81440 226500
rect 64380 226460 81440 226488
rect 64380 226448 64386 226460
rect 81434 226448 81440 226460
rect 81492 226448 81498 226500
rect 91462 226448 91468 226500
rect 91520 226488 91526 226500
rect 109678 226488 109684 226500
rect 91520 226460 109684 226488
rect 91520 226448 91526 226460
rect 109678 226448 109684 226460
rect 109736 226448 109742 226500
rect 119430 226448 119436 226500
rect 119488 226488 119494 226500
rect 137646 226488 137652 226500
rect 119488 226460 137652 226488
rect 119488 226448 119494 226460
rect 137646 226448 137652 226460
rect 137704 226448 137710 226500
rect 156322 226448 156328 226500
rect 156380 226488 156386 226500
rect 178678 226488 178684 226500
rect 156380 226460 178684 226488
rect 156380 226448 156386 226460
rect 178678 226448 178684 226460
rect 178736 226448 178742 226500
rect 232498 226448 232504 226500
rect 232556 226488 232562 226500
rect 249702 226488 249708 226500
rect 232556 226460 249708 226488
rect 232556 226448 232562 226460
rect 249702 226448 249708 226460
rect 249760 226448 249766 226500
rect 260190 226448 260196 226500
rect 260248 226488 260254 226500
rect 277670 226488 277676 226500
rect 260248 226460 277676 226488
rect 260248 226448 260254 226460
rect 277670 226448 277676 226460
rect 277728 226448 277734 226500
rect 287514 226448 287520 226500
rect 287572 226488 287578 226500
rect 305362 226488 305368 226500
rect 287572 226460 305368 226488
rect 287572 226448 287578 226460
rect 305362 226448 305368 226460
rect 305420 226448 305426 226500
rect 345658 226448 345664 226500
rect 345716 226488 345722 226500
rect 361666 226488 361672 226500
rect 345716 226460 361672 226488
rect 345716 226448 345722 226460
rect 361666 226448 361672 226460
rect 361724 226448 361730 226500
rect 371510 226448 371516 226500
rect 371568 226488 371574 226500
rect 389358 226488 389364 226500
rect 371568 226460 389364 226488
rect 371568 226448 371574 226460
rect 389358 226448 389364 226460
rect 389416 226448 389422 226500
rect 399478 226448 399484 226500
rect 399536 226488 399542 226500
rect 417694 226488 417700 226500
rect 399536 226460 417700 226488
rect 399536 226448 399542 226460
rect 417694 226448 417700 226460
rect 417752 226448 417758 226500
rect 456150 226448 456156 226500
rect 456208 226488 456214 226500
rect 473354 226488 473360 226500
rect 456208 226460 473360 226488
rect 456208 226448 456214 226460
rect 473354 226448 473360 226460
rect 473412 226448 473418 226500
rect 483474 226448 483480 226500
rect 483532 226488 483538 226500
rect 501690 226488 501696 226500
rect 483532 226460 501696 226488
rect 483532 226448 483538 226460
rect 501690 226448 501696 226460
rect 501748 226448 501754 226500
rect 36906 226380 36912 226432
rect 36964 226420 36970 226432
rect 63310 226420 63316 226432
rect 36964 226392 63316 226420
rect 36964 226380 36970 226392
rect 63310 226380 63316 226392
rect 63368 226380 63374 226432
rect 66898 226380 66904 226432
rect 66956 226420 66962 226432
rect 91094 226420 91100 226432
rect 66956 226392 91100 226420
rect 66956 226380 66962 226392
rect 91094 226380 91100 226392
rect 91152 226380 91158 226432
rect 94498 226380 94504 226432
rect 94556 226420 94562 226432
rect 119338 226420 119344 226432
rect 94556 226392 119344 226420
rect 94556 226380 94562 226392
rect 119338 226380 119344 226392
rect 119396 226380 119402 226432
rect 120718 226380 120724 226432
rect 120776 226420 120782 226432
rect 147306 226420 147312 226432
rect 120776 226392 147312 226420
rect 120776 226380 120782 226392
rect 147306 226380 147312 226392
rect 147364 226380 147370 226432
rect 148410 226380 148416 226432
rect 148468 226420 148474 226432
rect 175366 226420 175372 226432
rect 148468 226392 175372 226420
rect 148468 226380 148474 226392
rect 175366 226380 175372 226392
rect 175424 226380 175430 226432
rect 177298 226380 177304 226432
rect 177356 226420 177362 226432
rect 203334 226420 203340 226432
rect 177356 226392 203340 226420
rect 177356 226380 177362 226392
rect 203334 226380 203340 226392
rect 203392 226380 203398 226432
rect 204898 226380 204904 226432
rect 204956 226420 204962 226432
rect 231026 226420 231032 226432
rect 204956 226392 231032 226420
rect 204956 226380 204962 226392
rect 231026 226380 231032 226392
rect 231084 226380 231090 226432
rect 232590 226380 232596 226432
rect 232648 226420 232654 226432
rect 259362 226420 259368 226432
rect 232648 226392 259368 226420
rect 232648 226380 232654 226392
rect 259362 226380 259368 226392
rect 259420 226380 259426 226432
rect 268010 226380 268016 226432
rect 268068 226420 268074 226432
rect 287698 226420 287704 226432
rect 268068 226392 287704 226420
rect 268068 226380 268074 226392
rect 287698 226380 287704 226392
rect 287756 226380 287762 226432
rect 315482 226380 315488 226432
rect 315540 226420 315546 226432
rect 333698 226420 333704 226432
rect 315540 226392 333704 226420
rect 315540 226380 315546 226392
rect 333698 226380 333704 226392
rect 333756 226380 333762 226432
rect 352006 226380 352012 226432
rect 352064 226420 352070 226432
rect 374638 226420 374644 226432
rect 352064 226392 374644 226420
rect 352064 226380 352070 226392
rect 374638 226380 374644 226392
rect 374696 226380 374702 226432
rect 428550 226380 428556 226432
rect 428608 226420 428614 226432
rect 445662 226420 445668 226432
rect 428608 226392 445668 226420
rect 428608 226380 428614 226392
rect 445662 226380 445668 226392
rect 445720 226380 445726 226432
rect 464338 226380 464344 226432
rect 464396 226420 464402 226432
rect 483658 226420 483664 226432
rect 464396 226392 483664 226420
rect 464396 226380 464402 226392
rect 483658 226380 483664 226392
rect 483716 226380 483722 226432
rect 511442 226380 511448 226432
rect 511500 226420 511506 226432
rect 529658 226420 529664 226432
rect 511500 226392 529664 226420
rect 511500 226380 511506 226392
rect 529658 226380 529664 226392
rect 529716 226380 529722 226432
rect 542998 226380 543004 226432
rect 543056 226420 543062 226432
rect 557534 226420 557540 226432
rect 543056 226392 557540 226420
rect 543056 226380 543062 226392
rect 557534 226380 557540 226392
rect 557592 226380 557598 226432
rect 212350 226312 212356 226364
rect 212408 226352 212414 226364
rect 232682 226352 232688 226364
rect 212408 226324 232688 226352
rect 212408 226312 212414 226324
rect 232682 226312 232688 226324
rect 232740 226312 232746 226364
rect 260098 226312 260104 226364
rect 260156 226352 260162 226364
rect 287330 226352 287336 226364
rect 260156 226324 287336 226352
rect 260156 226312 260162 226324
rect 287330 226312 287336 226324
rect 287388 226312 287394 226364
rect 289078 226312 289084 226364
rect 289136 226352 289142 226364
rect 315022 226352 315028 226364
rect 289136 226324 315028 226352
rect 289136 226312 289142 226324
rect 315022 226312 315028 226324
rect 315080 226312 315086 226364
rect 316678 226312 316684 226364
rect 316736 226352 316742 226364
rect 343358 226352 343364 226364
rect 316736 226324 343364 226352
rect 316736 226312 316742 226324
rect 343358 226312 343364 226324
rect 343416 226312 343422 226364
rect 344278 226312 344284 226364
rect 344336 226352 344342 226364
rect 371326 226352 371332 226364
rect 344336 226324 371332 226352
rect 344336 226312 344342 226324
rect 371326 226312 371332 226324
rect 371384 226312 371390 226364
rect 373258 226312 373264 226364
rect 373316 226352 373322 226364
rect 399018 226352 399024 226364
rect 373316 226324 399024 226352
rect 373316 226312 373322 226324
rect 399018 226312 399024 226324
rect 399076 226312 399082 226364
rect 400858 226312 400864 226364
rect 400916 226352 400922 226364
rect 427354 226352 427360 226364
rect 400916 226324 427360 226352
rect 400916 226312 400922 226324
rect 427354 226312 427360 226324
rect 427412 226312 427418 226364
rect 428458 226312 428464 226364
rect 428516 226352 428522 226364
rect 455322 226352 455328 226364
rect 428516 226324 455328 226352
rect 428516 226312 428522 226324
rect 455322 226312 455328 226324
rect 455380 226312 455386 226364
rect 456058 226312 456064 226364
rect 456116 226352 456122 226364
rect 483014 226352 483020 226364
rect 456116 226324 483020 226352
rect 456116 226312 456122 226324
rect 483014 226312 483020 226324
rect 483072 226312 483078 226364
rect 485038 226312 485044 226364
rect 485096 226352 485102 226364
rect 511350 226352 511356 226364
rect 485096 226324 511356 226352
rect 485096 226312 485102 226324
rect 511350 226312 511356 226324
rect 511408 226312 511414 226364
rect 512638 226312 512644 226364
rect 512696 226352 512702 226364
rect 539318 226352 539324 226364
rect 512696 226324 539324 226352
rect 512696 226312 512702 226324
rect 539318 226312 539324 226324
rect 539376 226312 539382 226364
rect 540238 226312 540244 226364
rect 540296 226352 540302 226364
rect 567194 226352 567200 226364
rect 540296 226324 567200 226352
rect 540296 226312 540302 226324
rect 567194 226312 567200 226324
rect 567252 226312 567258 226364
rect 37918 225564 37924 225616
rect 37976 225604 37982 225616
rect 545758 225604 545764 225616
rect 37976 225576 545764 225604
rect 37976 225564 37982 225576
rect 545758 225564 545764 225576
rect 545816 225564 545822 225616
rect 35618 223592 35624 223644
rect 35676 223632 35682 223644
rect 36814 223632 36820 223644
rect 35676 223604 36820 223632
rect 35676 223592 35682 223604
rect 36814 223592 36820 223604
rect 36872 223592 36878 223644
rect 232682 207748 232688 207800
rect 232740 207788 232746 207800
rect 239766 207788 239772 207800
rect 232740 207760 239772 207788
rect 232740 207748 232746 207760
rect 239766 207748 239772 207760
rect 239824 207748 239830 207800
rect 428642 207612 428648 207664
rect 428700 207652 428706 207664
rect 435726 207652 435732 207664
rect 428700 207624 435732 207652
rect 428700 207612 428706 207624
rect 435726 207612 435732 207624
rect 435784 207612 435790 207664
rect 483658 207408 483664 207460
rect 483716 207448 483722 207460
rect 491662 207448 491668 207460
rect 483716 207420 491668 207448
rect 483716 207408 483722 207420
rect 491662 207408 491668 207420
rect 491720 207408 491726 207460
rect 63586 207340 63592 207392
rect 63644 207380 63650 207392
rect 64322 207380 64328 207392
rect 63644 207352 64328 207380
rect 63644 207340 63650 207352
rect 64322 207340 64328 207352
rect 64380 207340 64386 207392
rect 259730 207340 259736 207392
rect 259788 207380 259794 207392
rect 260190 207380 260196 207392
rect 259788 207352 260196 207380
rect 259788 207340 259794 207352
rect 260190 207340 260196 207352
rect 260248 207340 260254 207392
rect 316770 207340 316776 207392
rect 316828 207380 316834 207392
rect 323670 207380 323676 207392
rect 316828 207352 323676 207380
rect 316828 207340 316834 207352
rect 323670 207340 323676 207352
rect 323728 207340 323734 207392
rect 455690 207340 455696 207392
rect 455748 207380 455754 207392
rect 456150 207380 456156 207392
rect 455748 207352 456156 207380
rect 455748 207340 455754 207352
rect 456150 207340 456156 207352
rect 456208 207340 456214 207392
rect 512730 207272 512736 207324
rect 512788 207312 512794 207324
rect 519630 207312 519636 207324
rect 512788 207284 519636 207312
rect 512788 207272 512794 207284
rect 519630 207272 519636 207284
rect 519688 207272 519694 207324
rect 287698 207136 287704 207188
rect 287756 207176 287762 207188
rect 295702 207176 295708 207188
rect 287756 207148 295708 207176
rect 287756 207136 287762 207148
rect 295702 207136 295708 207148
rect 295760 207136 295766 207188
rect 13722 205572 13728 205624
rect 13780 205612 13786 205624
rect 66254 205612 66260 205624
rect 13780 205584 66260 205612
rect 13780 205572 13786 205584
rect 66254 205572 66260 205584
rect 66312 205572 66318 205624
rect 70302 205572 70308 205624
rect 70360 205612 70366 205624
rect 121454 205612 121460 205624
rect 70360 205584 121460 205612
rect 70360 205572 70366 205584
rect 121454 205572 121460 205584
rect 121512 205572 121518 205624
rect 126882 205572 126888 205624
rect 126940 205612 126946 205624
rect 178034 205612 178040 205624
rect 126940 205584 178040 205612
rect 126940 205572 126946 205584
rect 178034 205572 178040 205584
rect 178092 205572 178098 205624
rect 209682 205572 209688 205624
rect 209740 205612 209746 205624
rect 262214 205612 262220 205624
rect 209740 205584 262220 205612
rect 209740 205572 209746 205584
rect 262214 205572 262220 205584
rect 262272 205572 262278 205624
rect 266262 205572 266268 205624
rect 266320 205612 266326 205624
rect 317414 205612 317420 205624
rect 266320 205584 317420 205612
rect 266320 205572 266326 205584
rect 317414 205572 317420 205584
rect 317472 205572 317478 205624
rect 322842 205572 322848 205624
rect 322900 205612 322906 205624
rect 373994 205612 374000 205624
rect 322900 205584 374000 205612
rect 322900 205572 322906 205584
rect 373994 205572 374000 205584
rect 374052 205572 374058 205624
rect 405642 205572 405648 205624
rect 405700 205612 405706 205624
rect 458174 205612 458180 205624
rect 405700 205584 458180 205612
rect 405700 205572 405706 205584
rect 458174 205572 458180 205584
rect 458232 205572 458238 205624
rect 489822 205572 489828 205624
rect 489880 205612 489886 205624
rect 542354 205612 542360 205624
rect 489880 205584 542360 205612
rect 489880 205572 489886 205584
rect 542354 205572 542360 205584
rect 542412 205572 542418 205624
rect 35618 205504 35624 205556
rect 35676 205544 35682 205556
rect 36998 205544 37004 205556
rect 35676 205516 37004 205544
rect 35676 205504 35682 205516
rect 36998 205504 37004 205516
rect 37056 205504 37062 205556
rect 42702 205504 42708 205556
rect 42760 205544 42766 205556
rect 93854 205544 93860 205556
rect 42760 205516 93860 205544
rect 42760 205504 42766 205516
rect 93854 205504 93860 205516
rect 93912 205504 93918 205556
rect 97902 205504 97908 205556
rect 97960 205544 97966 205556
rect 149054 205544 149060 205556
rect 97960 205516 149060 205544
rect 97960 205504 97966 205516
rect 149054 205504 149060 205516
rect 149112 205504 149118 205556
rect 154482 205504 154488 205556
rect 154540 205544 154546 205556
rect 205634 205544 205640 205556
rect 154540 205516 205640 205544
rect 154540 205504 154546 205516
rect 205634 205504 205640 205516
rect 205692 205504 205698 205556
rect 238662 205504 238668 205556
rect 238720 205544 238726 205556
rect 289814 205544 289820 205556
rect 238720 205516 289820 205544
rect 238720 205504 238726 205516
rect 289814 205504 289820 205516
rect 289872 205504 289878 205556
rect 293862 205504 293868 205556
rect 293920 205544 293926 205556
rect 345014 205544 345020 205556
rect 293920 205516 345020 205544
rect 293920 205504 293926 205516
rect 345014 205504 345020 205516
rect 345072 205504 345078 205556
rect 350442 205504 350448 205556
rect 350500 205544 350506 205556
rect 401594 205544 401600 205556
rect 350500 205516 401600 205544
rect 350500 205504 350506 205516
rect 401594 205504 401600 205516
rect 401652 205504 401658 205556
rect 427722 205504 427728 205556
rect 427780 205544 427786 205556
rect 428550 205544 428556 205556
rect 427780 205516 428556 205544
rect 427780 205504 427786 205516
rect 428550 205504 428556 205516
rect 428608 205504 428614 205556
rect 434622 205504 434628 205556
rect 434680 205544 434686 205556
rect 485774 205544 485780 205556
rect 434680 205516 485780 205544
rect 434680 205504 434686 205516
rect 485774 205504 485780 205516
rect 485832 205504 485838 205556
rect 518802 205504 518808 205556
rect 518860 205544 518866 205556
rect 569954 205544 569960 205556
rect 518860 205516 569960 205544
rect 518860 205504 518866 205516
rect 569954 205504 569960 205516
rect 570012 205504 570018 205556
rect 182082 205436 182088 205488
rect 182140 205476 182146 205488
rect 233234 205476 233240 205488
rect 182140 205448 233240 205476
rect 182140 205436 182146 205448
rect 233234 205436 233240 205448
rect 233292 205436 233298 205488
rect 343634 205436 343640 205488
rect 343692 205476 343698 205488
rect 345658 205476 345664 205488
rect 343692 205448 345664 205476
rect 343692 205436 343698 205448
rect 345658 205436 345664 205448
rect 345716 205436 345722 205488
rect 378042 205436 378048 205488
rect 378100 205476 378106 205488
rect 429194 205476 429200 205488
rect 378100 205448 429200 205476
rect 378100 205436 378106 205448
rect 429194 205436 429200 205448
rect 429252 205436 429258 205488
rect 462222 205436 462228 205488
rect 462280 205476 462286 205488
rect 513374 205476 513380 205488
rect 462280 205448 513380 205476
rect 462280 205436 462286 205448
rect 513374 205436 513380 205448
rect 513432 205436 513438 205488
rect 539502 205436 539508 205488
rect 539560 205476 539566 205488
rect 542998 205476 543004 205488
rect 539560 205448 543004 205476
rect 539560 205436 539566 205448
rect 542998 205436 543004 205448
rect 543056 205436 543062 205488
rect 178678 202784 178684 202836
rect 178736 202824 178742 202836
rect 184014 202824 184020 202836
rect 178736 202796 184020 202824
rect 178736 202784 178742 202796
rect 184014 202784 184020 202796
rect 184072 202784 184078 202836
rect 374638 202784 374644 202836
rect 374696 202824 374702 202836
rect 379698 202824 379704 202836
rect 374696 202796 379704 202824
rect 374696 202784 374702 202796
rect 379698 202784 379704 202796
rect 379756 202784 379762 202836
rect 15194 202716 15200 202768
rect 15252 202756 15258 202768
rect 43622 202756 43628 202768
rect 15252 202728 43628 202756
rect 15252 202716 15258 202728
rect 43622 202716 43628 202728
rect 43680 202716 43686 202768
rect 69658 202716 69664 202768
rect 69716 202756 69722 202768
rect 567194 202756 567200 202768
rect 69716 202728 567200 202756
rect 69716 202716 69722 202728
rect 567194 202716 567200 202728
rect 567252 202716 567258 202768
rect 25682 202648 25688 202700
rect 25740 202688 25746 202700
rect 36906 202688 36912 202700
rect 25740 202660 36912 202688
rect 25740 202648 25746 202660
rect 36906 202648 36912 202660
rect 36964 202648 36970 202700
rect 53558 202648 53564 202700
rect 53616 202688 53622 202700
rect 66898 202688 66904 202700
rect 53616 202660 66904 202688
rect 53616 202648 53622 202660
rect 66898 202648 66904 202660
rect 66956 202648 66962 202700
rect 71866 202648 71872 202700
rect 71924 202688 71930 202700
rect 100018 202688 100024 202700
rect 71924 202660 100024 202688
rect 71924 202648 71930 202660
rect 100018 202648 100024 202660
rect 100076 202648 100082 202700
rect 127710 202688 127716 202700
rect 103486 202660 127716 202688
rect 42886 202580 42892 202632
rect 42944 202620 42950 202632
rect 72050 202620 72056 202632
rect 42944 202592 72056 202620
rect 42944 202580 42950 202592
rect 72050 202580 72056 202592
rect 72108 202580 72114 202632
rect 81986 202580 81992 202632
rect 82044 202620 82050 202632
rect 94498 202620 94504 202632
rect 82044 202592 94504 202620
rect 82044 202580 82050 202592
rect 94498 202580 94504 202592
rect 94556 202580 94562 202632
rect 99466 202580 99472 202632
rect 99524 202620 99530 202632
rect 103486 202620 103514 202660
rect 127710 202648 127716 202660
rect 127768 202648 127774 202700
rect 156046 202688 156052 202700
rect 132466 202660 156052 202688
rect 99524 202592 103514 202620
rect 99524 202580 99530 202592
rect 109678 202580 109684 202632
rect 109736 202620 109742 202632
rect 120718 202620 120724 202632
rect 109736 202592 120724 202620
rect 109736 202580 109742 202592
rect 120718 202580 120724 202592
rect 120776 202580 120782 202632
rect 127066 202580 127072 202632
rect 127124 202620 127130 202632
rect 132466 202620 132494 202660
rect 156046 202648 156052 202660
rect 156104 202648 156110 202700
rect 165982 202648 165988 202700
rect 166040 202688 166046 202700
rect 177298 202688 177304 202700
rect 166040 202660 177304 202688
rect 166040 202648 166046 202660
rect 177298 202648 177304 202660
rect 177356 202648 177362 202700
rect 183646 202648 183652 202700
rect 183704 202688 183710 202700
rect 211706 202688 211712 202700
rect 183704 202660 211712 202688
rect 183704 202648 183710 202660
rect 211706 202648 211712 202660
rect 211764 202648 211770 202700
rect 222010 202648 222016 202700
rect 222068 202688 222074 202700
rect 232590 202688 232596 202700
rect 222068 202660 232596 202688
rect 222068 202648 222074 202660
rect 232590 202648 232596 202660
rect 232648 202648 232654 202700
rect 238846 202648 238852 202700
rect 238904 202688 238910 202700
rect 268010 202688 268016 202700
rect 238904 202660 268016 202688
rect 238904 202648 238910 202660
rect 268010 202648 268016 202660
rect 268068 202648 268074 202700
rect 277670 202648 277676 202700
rect 277728 202688 277734 202700
rect 289078 202688 289084 202700
rect 277728 202660 289084 202688
rect 277728 202648 277734 202660
rect 289078 202648 289084 202660
rect 289136 202648 289142 202700
rect 306006 202648 306012 202700
rect 306064 202688 306070 202700
rect 316678 202688 316684 202700
rect 306064 202660 316684 202688
rect 306064 202648 306070 202660
rect 316678 202648 316684 202660
rect 316736 202648 316742 202700
rect 323026 202648 323032 202700
rect 323084 202688 323090 202700
rect 352006 202688 352012 202700
rect 323084 202660 352012 202688
rect 323084 202648 323090 202660
rect 352006 202648 352012 202660
rect 352064 202648 352070 202700
rect 361666 202648 361672 202700
rect 361724 202688 361730 202700
rect 373258 202688 373264 202700
rect 361724 202660 373264 202688
rect 361724 202648 361730 202660
rect 373258 202648 373264 202660
rect 373316 202648 373322 202700
rect 379606 202648 379612 202700
rect 379664 202688 379670 202700
rect 408034 202688 408040 202700
rect 379664 202660 408040 202688
rect 379664 202648 379670 202660
rect 408034 202648 408040 202660
rect 408092 202648 408098 202700
rect 417694 202648 417700 202700
rect 417752 202688 417758 202700
rect 428458 202688 428464 202700
rect 417752 202660 428464 202688
rect 417752 202648 417758 202660
rect 428458 202648 428464 202660
rect 428516 202648 428522 202700
rect 434806 202648 434812 202700
rect 434864 202688 434870 202700
rect 463694 202688 463700 202700
rect 434864 202660 463700 202688
rect 434864 202648 434870 202660
rect 463694 202648 463700 202660
rect 463752 202648 463758 202700
rect 473998 202648 474004 202700
rect 474056 202688 474062 202700
rect 485038 202688 485044 202700
rect 474056 202660 485044 202688
rect 474056 202648 474062 202660
rect 485038 202648 485044 202660
rect 485096 202648 485102 202700
rect 501690 202648 501696 202700
rect 501748 202688 501754 202700
rect 512638 202688 512644 202700
rect 501748 202660 512644 202688
rect 501748 202648 501754 202660
rect 512638 202648 512644 202660
rect 512696 202648 512702 202700
rect 518986 202648 518992 202700
rect 519044 202688 519050 202700
rect 547874 202688 547880 202700
rect 519044 202660 547880 202688
rect 519044 202648 519050 202660
rect 547874 202648 547880 202660
rect 547932 202648 547938 202700
rect 127124 202592 132494 202620
rect 127124 202580 127130 202592
rect 137922 202580 137928 202632
rect 137980 202620 137986 202632
rect 148410 202620 148416 202632
rect 137980 202592 148416 202620
rect 137980 202580 137986 202592
rect 148410 202580 148416 202592
rect 148468 202580 148474 202632
rect 193674 202580 193680 202632
rect 193732 202620 193738 202632
rect 204898 202620 204904 202632
rect 193732 202592 204904 202620
rect 193732 202580 193738 202592
rect 204898 202580 204904 202592
rect 204956 202580 204962 202632
rect 249518 202580 249524 202632
rect 249576 202620 249582 202632
rect 260098 202620 260104 202632
rect 249576 202592 260104 202620
rect 249576 202580 249582 202592
rect 260098 202580 260104 202592
rect 260156 202580 260162 202632
rect 333882 202580 333888 202632
rect 333940 202620 333946 202632
rect 344278 202620 344284 202632
rect 333940 202592 344284 202620
rect 333940 202580 333946 202592
rect 344278 202580 344284 202592
rect 344336 202580 344342 202632
rect 390002 202580 390008 202632
rect 390060 202620 390066 202632
rect 400858 202620 400864 202632
rect 390060 202592 400864 202620
rect 390060 202580 390066 202592
rect 400858 202580 400864 202592
rect 400916 202580 400922 202632
rect 445662 202580 445668 202632
rect 445720 202620 445726 202632
rect 456058 202620 456064 202632
rect 445720 202592 456064 202620
rect 445720 202580 445726 202592
rect 456058 202580 456064 202592
rect 456116 202580 456122 202632
rect 529658 202580 529664 202632
rect 529716 202620 529722 202632
rect 540238 202620 540244 202632
rect 529716 202592 540244 202620
rect 529716 202580 529722 202592
rect 540238 202580 540244 202592
rect 540296 202580 540302 202632
rect 36722 202512 36728 202564
rect 36780 202552 36786 202564
rect 557534 202552 557540 202564
rect 36780 202524 557540 202552
rect 36780 202512 36786 202524
rect 557534 202512 557540 202524
rect 557592 202512 557598 202564
rect 16022 200744 16028 200796
rect 16080 200784 16086 200796
rect 547874 200784 547880 200796
rect 16080 200756 547880 200784
rect 16080 200744 16086 200756
rect 547874 200744 547880 200756
rect 547932 200744 547938 200796
rect 25682 200336 25688 200388
rect 25740 200376 25746 200388
rect 71038 200376 71044 200388
rect 25740 200348 71044 200376
rect 25740 200336 25746 200348
rect 71038 200336 71044 200348
rect 71096 200336 71102 200388
rect 212258 200336 212264 200388
rect 212316 200376 212322 200388
rect 232682 200376 232688 200388
rect 212316 200348 232688 200376
rect 212316 200336 212322 200348
rect 232682 200336 232688 200348
rect 232740 200336 232746 200388
rect 296346 200336 296352 200388
rect 296404 200376 296410 200388
rect 316770 200376 316776 200388
rect 296404 200348 316776 200376
rect 296404 200336 296410 200348
rect 316770 200336 316776 200348
rect 316828 200336 316834 200388
rect 408034 200336 408040 200388
rect 408092 200376 408098 200388
rect 428642 200376 428648 200388
rect 408092 200348 428648 200376
rect 408092 200336 408098 200348
rect 428642 200336 428648 200348
rect 428700 200336 428706 200388
rect 492030 200336 492036 200388
rect 492088 200376 492094 200388
rect 512730 200376 512736 200388
rect 492088 200348 512736 200376
rect 492088 200336 492094 200348
rect 512730 200336 512736 200348
rect 512788 200336 512794 200388
rect 36906 200268 36912 200320
rect 36964 200308 36970 200320
rect 53650 200308 53656 200320
rect 36964 200280 53656 200308
rect 36964 200268 36970 200280
rect 53650 200268 53656 200280
rect 53708 200268 53714 200320
rect 148410 200268 148416 200320
rect 148468 200308 148474 200320
rect 165614 200308 165620 200320
rect 148468 200280 165620 200308
rect 148468 200268 148474 200280
rect 165614 200268 165620 200280
rect 165672 200268 165678 200320
rect 175458 200268 175464 200320
rect 175516 200308 175522 200320
rect 193674 200308 193680 200320
rect 175516 200280 193680 200308
rect 175516 200268 175522 200280
rect 193674 200268 193680 200280
rect 193732 200268 193738 200320
rect 203518 200268 203524 200320
rect 203576 200308 203582 200320
rect 221366 200308 221372 200320
rect 203576 200280 221372 200308
rect 203576 200268 203582 200280
rect 221366 200268 221372 200280
rect 221424 200268 221430 200320
rect 260190 200268 260196 200320
rect 260248 200308 260254 200320
rect 277670 200308 277676 200320
rect 260248 200280 277676 200308
rect 260248 200268 260254 200280
rect 277670 200268 277676 200280
rect 277728 200268 277734 200320
rect 287514 200268 287520 200320
rect 287572 200308 287578 200320
rect 305362 200308 305368 200320
rect 287572 200280 305368 200308
rect 287572 200268 287578 200280
rect 305362 200268 305368 200280
rect 305420 200268 305426 200320
rect 345658 200268 345664 200320
rect 345716 200308 345722 200320
rect 361666 200308 361672 200320
rect 345716 200280 361672 200308
rect 345716 200268 345722 200280
rect 361666 200268 361672 200280
rect 361724 200268 361730 200320
rect 371510 200268 371516 200320
rect 371568 200308 371574 200320
rect 389358 200308 389364 200320
rect 371568 200280 389364 200308
rect 371568 200268 371574 200280
rect 389358 200268 389364 200280
rect 389416 200268 389422 200320
rect 399478 200268 399484 200320
rect 399536 200308 399542 200320
rect 417694 200308 417700 200320
rect 399536 200280 417700 200308
rect 399536 200268 399542 200280
rect 417694 200268 417700 200280
rect 417752 200268 417758 200320
rect 456150 200268 456156 200320
rect 456208 200308 456214 200320
rect 473538 200308 473544 200320
rect 456208 200280 473544 200308
rect 456208 200268 456214 200280
rect 473538 200268 473544 200280
rect 473596 200268 473602 200320
rect 483474 200268 483480 200320
rect 483532 200308 483538 200320
rect 501690 200308 501696 200320
rect 483532 200280 501696 200308
rect 483532 200268 483538 200280
rect 501690 200268 501696 200280
rect 501748 200268 501754 200320
rect 36998 200200 37004 200252
rect 37056 200240 37062 200252
rect 63310 200240 63316 200252
rect 37056 200212 63316 200240
rect 37056 200200 37062 200212
rect 63310 200200 63316 200212
rect 63368 200200 63374 200252
rect 64322 200200 64328 200252
rect 64380 200240 64386 200252
rect 81434 200240 81440 200252
rect 64380 200212 81440 200240
rect 64380 200200 64386 200212
rect 81434 200200 81440 200212
rect 81492 200200 81498 200252
rect 91462 200200 91468 200252
rect 91520 200240 91526 200252
rect 109678 200240 109684 200252
rect 91520 200212 109684 200240
rect 91520 200200 91526 200212
rect 109678 200200 109684 200212
rect 109736 200200 109742 200252
rect 119430 200200 119436 200252
rect 119488 200240 119494 200252
rect 137646 200240 137652 200252
rect 119488 200212 137652 200240
rect 119488 200200 119494 200212
rect 137646 200200 137652 200212
rect 137704 200200 137710 200252
rect 156322 200200 156328 200252
rect 156380 200240 156386 200252
rect 178678 200240 178684 200252
rect 156380 200212 178684 200240
rect 156380 200200 156386 200212
rect 178678 200200 178684 200212
rect 178736 200200 178742 200252
rect 232590 200200 232596 200252
rect 232648 200240 232654 200252
rect 249702 200240 249708 200252
rect 232648 200212 249708 200240
rect 232648 200200 232654 200212
rect 249702 200200 249708 200212
rect 249760 200200 249766 200252
rect 268010 200200 268016 200252
rect 268068 200240 268074 200252
rect 287698 200240 287704 200252
rect 268068 200212 287704 200240
rect 268068 200200 268074 200212
rect 287698 200200 287704 200212
rect 287756 200200 287762 200252
rect 315482 200200 315488 200252
rect 315540 200240 315546 200252
rect 333698 200240 333704 200252
rect 315540 200212 333704 200240
rect 315540 200200 315546 200212
rect 333698 200200 333704 200212
rect 333756 200200 333762 200252
rect 352006 200200 352012 200252
rect 352064 200240 352070 200252
rect 374638 200240 374644 200252
rect 352064 200212 374644 200240
rect 352064 200200 352070 200212
rect 374638 200200 374644 200212
rect 374696 200200 374702 200252
rect 428458 200200 428464 200252
rect 428516 200240 428522 200252
rect 445662 200240 445668 200252
rect 428516 200212 445668 200240
rect 428516 200200 428522 200212
rect 445662 200200 445668 200212
rect 445720 200200 445726 200252
rect 464338 200200 464344 200252
rect 464396 200240 464402 200252
rect 483658 200240 483664 200252
rect 464396 200212 483664 200240
rect 464396 200200 464402 200212
rect 483658 200200 483664 200212
rect 483716 200200 483722 200252
rect 511442 200200 511448 200252
rect 511500 200240 511506 200252
rect 529658 200240 529664 200252
rect 511500 200212 529664 200240
rect 511500 200200 511506 200212
rect 529658 200200 529664 200212
rect 529716 200200 529722 200252
rect 542998 200200 543004 200252
rect 543056 200240 543062 200252
rect 557534 200240 557540 200252
rect 543056 200212 557540 200240
rect 543056 200200 543062 200212
rect 557534 200200 557540 200212
rect 557592 200200 557598 200252
rect 69658 200132 69664 200184
rect 69716 200172 69722 200184
rect 91094 200172 91100 200184
rect 69716 200144 91100 200172
rect 69716 200132 69722 200144
rect 91094 200132 91100 200144
rect 91152 200132 91158 200184
rect 94498 200132 94504 200184
rect 94556 200172 94562 200184
rect 119338 200172 119344 200184
rect 94556 200144 119344 200172
rect 94556 200132 94562 200144
rect 119338 200132 119344 200144
rect 119396 200132 119402 200184
rect 120718 200132 120724 200184
rect 120776 200172 120782 200184
rect 147306 200172 147312 200184
rect 120776 200144 147312 200172
rect 120776 200132 120782 200144
rect 147306 200132 147312 200144
rect 147364 200132 147370 200184
rect 148318 200132 148324 200184
rect 148376 200172 148382 200184
rect 175274 200172 175280 200184
rect 148376 200144 175280 200172
rect 148376 200132 148382 200144
rect 175274 200132 175280 200144
rect 175332 200132 175338 200184
rect 177298 200132 177304 200184
rect 177356 200172 177362 200184
rect 203334 200172 203340 200184
rect 177356 200144 203340 200172
rect 177356 200132 177362 200144
rect 203334 200132 203340 200144
rect 203392 200132 203398 200184
rect 204898 200132 204904 200184
rect 204956 200172 204962 200184
rect 231026 200172 231032 200184
rect 204956 200144 231032 200172
rect 204956 200132 204962 200144
rect 231026 200132 231032 200144
rect 231084 200132 231090 200184
rect 232498 200132 232504 200184
rect 232556 200172 232562 200184
rect 259362 200172 259368 200184
rect 232556 200144 259368 200172
rect 232556 200132 232562 200144
rect 259362 200132 259368 200144
rect 259420 200132 259426 200184
rect 260098 200132 260104 200184
rect 260156 200172 260162 200184
rect 287330 200172 287336 200184
rect 260156 200144 287336 200172
rect 260156 200132 260162 200144
rect 287330 200132 287336 200144
rect 287388 200132 287394 200184
rect 289078 200132 289084 200184
rect 289136 200172 289142 200184
rect 315022 200172 315028 200184
rect 289136 200144 315028 200172
rect 289136 200132 289142 200144
rect 315022 200132 315028 200144
rect 315080 200132 315086 200184
rect 316678 200132 316684 200184
rect 316736 200172 316742 200184
rect 343358 200172 343364 200184
rect 316736 200144 343364 200172
rect 316736 200132 316742 200144
rect 343358 200132 343364 200144
rect 343416 200132 343422 200184
rect 344278 200132 344284 200184
rect 344336 200172 344342 200184
rect 371326 200172 371332 200184
rect 344336 200144 371332 200172
rect 344336 200132 344342 200144
rect 371326 200132 371332 200144
rect 371384 200132 371390 200184
rect 373258 200132 373264 200184
rect 373316 200172 373322 200184
rect 399018 200172 399024 200184
rect 373316 200144 399024 200172
rect 373316 200132 373322 200144
rect 399018 200132 399024 200144
rect 399076 200132 399082 200184
rect 400858 200132 400864 200184
rect 400916 200172 400922 200184
rect 427354 200172 427360 200184
rect 400916 200144 427360 200172
rect 400916 200132 400922 200144
rect 427354 200132 427360 200144
rect 427412 200132 427418 200184
rect 428550 200132 428556 200184
rect 428608 200172 428614 200184
rect 455322 200172 455328 200184
rect 428608 200144 455328 200172
rect 428608 200132 428614 200144
rect 455322 200132 455328 200144
rect 455380 200132 455386 200184
rect 456058 200132 456064 200184
rect 456116 200172 456122 200184
rect 483198 200172 483204 200184
rect 456116 200144 483204 200172
rect 456116 200132 456122 200144
rect 483198 200132 483204 200144
rect 483256 200132 483262 200184
rect 485038 200132 485044 200184
rect 485096 200172 485102 200184
rect 511350 200172 511356 200184
rect 485096 200144 511356 200172
rect 485096 200132 485102 200144
rect 511350 200132 511356 200144
rect 511408 200132 511414 200184
rect 512638 200132 512644 200184
rect 512696 200172 512702 200184
rect 539318 200172 539324 200184
rect 512696 200144 539324 200172
rect 512696 200132 512702 200144
rect 539318 200132 539324 200144
rect 539376 200132 539382 200184
rect 540238 200132 540244 200184
rect 540296 200172 540302 200184
rect 567194 200172 567200 200184
rect 540296 200144 567200 200172
rect 540296 200132 540302 200144
rect 567194 200132 567200 200144
rect 567252 200132 567258 200184
rect 37918 197956 37924 198008
rect 37976 197996 37982 198008
rect 545758 197996 545764 198008
rect 37976 197968 545764 197996
rect 37976 197956 37982 197968
rect 545758 197956 545764 197968
rect 545816 197956 545822 198008
rect 35618 197344 35624 197396
rect 35676 197384 35682 197396
rect 36722 197384 36728 197396
rect 35676 197356 36728 197384
rect 35676 197344 35682 197356
rect 36722 197344 36728 197356
rect 36780 197344 36786 197396
rect 2958 187688 2964 187740
rect 3016 187728 3022 187740
rect 13170 187728 13176 187740
rect 3016 187700 13176 187728
rect 3016 187688 3022 187700
rect 13170 187688 13176 187700
rect 13228 187688 13234 187740
rect 63586 185580 63592 185632
rect 63644 185620 63650 185632
rect 64322 185620 64328 185632
rect 63644 185592 64328 185620
rect 63644 185580 63650 185592
rect 64322 185580 64328 185592
rect 64380 185580 64386 185632
rect 147674 185580 147680 185632
rect 147732 185620 147738 185632
rect 148410 185620 148416 185632
rect 147732 185592 148416 185620
rect 147732 185580 147738 185592
rect 148410 185580 148416 185592
rect 148468 185580 148474 185632
rect 259730 185580 259736 185632
rect 259788 185620 259794 185632
rect 260190 185620 260196 185632
rect 259788 185592 260196 185620
rect 259788 185580 259794 185592
rect 260190 185580 260196 185592
rect 260248 185580 260254 185632
rect 455690 185580 455696 185632
rect 455748 185620 455754 185632
rect 456150 185620 456156 185632
rect 455748 185592 456156 185620
rect 455748 185580 455754 185592
rect 456150 185580 456156 185592
rect 456208 185580 456214 185632
rect 428642 180072 428648 180124
rect 428700 180112 428706 180124
rect 435726 180112 435732 180124
rect 428700 180084 435732 180112
rect 428700 180072 428706 180084
rect 435726 180072 435732 180084
rect 435784 180072 435790 180124
rect 232682 179868 232688 179920
rect 232740 179908 232746 179920
rect 239766 179908 239772 179920
rect 232740 179880 239772 179908
rect 232740 179868 232746 179880
rect 239766 179868 239772 179880
rect 239824 179868 239830 179920
rect 512730 179800 512736 179852
rect 512788 179840 512794 179852
rect 519630 179840 519636 179852
rect 512788 179812 519636 179840
rect 512788 179800 512794 179812
rect 519630 179800 519636 179812
rect 519688 179800 519694 179852
rect 483658 179664 483664 179716
rect 483716 179704 483722 179716
rect 491662 179704 491668 179716
rect 483716 179676 491668 179704
rect 483716 179664 483722 179676
rect 491662 179664 491668 179676
rect 491720 179664 491726 179716
rect 287698 179392 287704 179444
rect 287756 179432 287762 179444
rect 295702 179432 295708 179444
rect 287756 179404 295708 179432
rect 287756 179392 287762 179404
rect 295702 179392 295708 179404
rect 295760 179392 295766 179444
rect 316770 179392 316776 179444
rect 316828 179432 316834 179444
rect 323670 179432 323676 179444
rect 316828 179404 323676 179432
rect 316828 179392 316834 179404
rect 323670 179392 323676 179404
rect 323728 179392 323734 179444
rect 13722 179324 13728 179376
rect 13780 179364 13786 179376
rect 66254 179364 66260 179376
rect 13780 179336 66260 179364
rect 13780 179324 13786 179336
rect 66254 179324 66260 179336
rect 66312 179324 66318 179376
rect 70302 179324 70308 179376
rect 70360 179364 70366 179376
rect 121454 179364 121460 179376
rect 70360 179336 121460 179364
rect 70360 179324 70366 179336
rect 121454 179324 121460 179336
rect 121512 179324 121518 179376
rect 126882 179324 126888 179376
rect 126940 179364 126946 179376
rect 178034 179364 178040 179376
rect 126940 179336 178040 179364
rect 126940 179324 126946 179336
rect 178034 179324 178040 179336
rect 178092 179324 178098 179376
rect 209682 179324 209688 179376
rect 209740 179364 209746 179376
rect 262214 179364 262220 179376
rect 209740 179336 262220 179364
rect 209740 179324 209746 179336
rect 262214 179324 262220 179336
rect 262272 179324 262278 179376
rect 266262 179324 266268 179376
rect 266320 179364 266326 179376
rect 317414 179364 317420 179376
rect 266320 179336 317420 179364
rect 266320 179324 266326 179336
rect 317414 179324 317420 179336
rect 317472 179324 317478 179376
rect 322842 179324 322848 179376
rect 322900 179364 322906 179376
rect 373994 179364 374000 179376
rect 322900 179336 374000 179364
rect 322900 179324 322906 179336
rect 373994 179324 374000 179336
rect 374052 179324 374058 179376
rect 405642 179324 405648 179376
rect 405700 179364 405706 179376
rect 458174 179364 458180 179376
rect 405700 179336 458180 179364
rect 405700 179324 405706 179336
rect 458174 179324 458180 179336
rect 458232 179324 458238 179376
rect 489822 179324 489828 179376
rect 489880 179364 489886 179376
rect 542354 179364 542360 179376
rect 489880 179336 542360 179364
rect 489880 179324 489886 179336
rect 542354 179324 542360 179336
rect 542412 179324 542418 179376
rect 35618 179256 35624 179308
rect 35676 179296 35682 179308
rect 36906 179296 36912 179308
rect 35676 179268 36912 179296
rect 35676 179256 35682 179268
rect 36906 179256 36912 179268
rect 36964 179256 36970 179308
rect 42702 179256 42708 179308
rect 42760 179296 42766 179308
rect 93854 179296 93860 179308
rect 42760 179268 93860 179296
rect 42760 179256 42766 179268
rect 93854 179256 93860 179268
rect 93912 179256 93918 179308
rect 97902 179256 97908 179308
rect 97960 179296 97966 179308
rect 149054 179296 149060 179308
rect 97960 179268 149060 179296
rect 97960 179256 97966 179268
rect 149054 179256 149060 179268
rect 149112 179256 149118 179308
rect 154482 179256 154488 179308
rect 154540 179296 154546 179308
rect 205634 179296 205640 179308
rect 154540 179268 205640 179296
rect 154540 179256 154546 179268
rect 205634 179256 205640 179268
rect 205692 179256 205698 179308
rect 231670 179256 231676 179308
rect 231728 179296 231734 179308
rect 232590 179296 232596 179308
rect 231728 179268 232596 179296
rect 231728 179256 231734 179268
rect 232590 179256 232596 179268
rect 232648 179256 232654 179308
rect 238662 179256 238668 179308
rect 238720 179296 238726 179308
rect 289814 179296 289820 179308
rect 238720 179268 289820 179296
rect 238720 179256 238726 179268
rect 289814 179256 289820 179268
rect 289872 179256 289878 179308
rect 293862 179256 293868 179308
rect 293920 179296 293926 179308
rect 293920 179268 335354 179296
rect 293920 179256 293926 179268
rect 182082 179188 182088 179240
rect 182140 179228 182146 179240
rect 233234 179228 233240 179240
rect 182140 179200 233240 179228
rect 182140 179188 182146 179200
rect 233234 179188 233240 179200
rect 233292 179188 233298 179240
rect 335326 179228 335354 179268
rect 343542 179256 343548 179308
rect 343600 179296 343606 179308
rect 345658 179296 345664 179308
rect 343600 179268 345664 179296
rect 343600 179256 343606 179268
rect 345658 179256 345664 179268
rect 345716 179256 345722 179308
rect 350442 179256 350448 179308
rect 350500 179296 350506 179308
rect 401594 179296 401600 179308
rect 350500 179268 401600 179296
rect 350500 179256 350506 179268
rect 401594 179256 401600 179268
rect 401652 179256 401658 179308
rect 434622 179256 434628 179308
rect 434680 179296 434686 179308
rect 485774 179296 485780 179308
rect 434680 179268 485780 179296
rect 434680 179256 434686 179268
rect 485774 179256 485780 179268
rect 485832 179256 485838 179308
rect 518802 179256 518808 179308
rect 518860 179296 518866 179308
rect 569954 179296 569960 179308
rect 518860 179268 569960 179296
rect 518860 179256 518866 179268
rect 569954 179256 569960 179268
rect 570012 179256 570018 179308
rect 345014 179228 345020 179240
rect 335326 179200 345020 179228
rect 345014 179188 345020 179200
rect 345072 179188 345078 179240
rect 378042 179188 378048 179240
rect 378100 179228 378106 179240
rect 429194 179228 429200 179240
rect 378100 179200 429200 179228
rect 378100 179188 378106 179200
rect 429194 179188 429200 179200
rect 429252 179188 429258 179240
rect 462222 179188 462228 179240
rect 462280 179228 462286 179240
rect 513374 179228 513380 179240
rect 462280 179200 513380 179228
rect 462280 179188 462286 179200
rect 513374 179188 513380 179200
rect 513432 179188 513438 179240
rect 42886 176604 42892 176656
rect 42944 176644 42950 176656
rect 72050 176644 72056 176656
rect 42944 176616 45554 176644
rect 42944 176604 42950 176616
rect 15194 176536 15200 176588
rect 15252 176576 15258 176588
rect 43990 176576 43996 176588
rect 15252 176548 43996 176576
rect 15252 176536 15258 176548
rect 43990 176536 43996 176548
rect 44048 176536 44054 176588
rect 45526 176576 45554 176616
rect 64846 176616 72056 176644
rect 64846 176576 64874 176616
rect 72050 176604 72056 176616
rect 72108 176604 72114 176656
rect 99466 176604 99472 176656
rect 99524 176644 99530 176656
rect 99524 176616 103514 176644
rect 99524 176604 99530 176616
rect 45526 176548 64874 176576
rect 71866 176536 71872 176588
rect 71924 176576 71930 176588
rect 100018 176576 100024 176588
rect 71924 176548 100024 176576
rect 71924 176536 71930 176548
rect 100018 176536 100024 176548
rect 100076 176536 100082 176588
rect 103486 176576 103514 176616
rect 127066 176604 127072 176656
rect 127124 176644 127130 176656
rect 127124 176616 132494 176644
rect 127124 176604 127130 176616
rect 127986 176576 127992 176588
rect 103486 176548 127992 176576
rect 127986 176536 127992 176548
rect 128044 176536 128050 176588
rect 132466 176576 132494 176616
rect 183646 176604 183652 176656
rect 183704 176644 183710 176656
rect 183704 176616 190454 176644
rect 183704 176604 183710 176616
rect 156046 176576 156052 176588
rect 132466 176548 156052 176576
rect 156046 176536 156052 176548
rect 156104 176536 156110 176588
rect 165982 176536 165988 176588
rect 166040 176576 166046 176588
rect 177298 176576 177304 176588
rect 166040 176548 177304 176576
rect 166040 176536 166046 176548
rect 177298 176536 177304 176548
rect 177356 176536 177362 176588
rect 178678 176536 178684 176588
rect 178736 176576 178742 176588
rect 184014 176576 184020 176588
rect 178736 176548 184020 176576
rect 178736 176536 178742 176548
rect 184014 176536 184020 176548
rect 184072 176536 184078 176588
rect 190426 176576 190454 176616
rect 374638 176604 374644 176656
rect 374696 176644 374702 176656
rect 379698 176644 379704 176656
rect 374696 176616 379704 176644
rect 374696 176604 374702 176616
rect 379698 176604 379704 176616
rect 379756 176604 379762 176656
rect 539318 176604 539324 176656
rect 539376 176644 539382 176656
rect 542998 176644 543004 176656
rect 539376 176616 543004 176644
rect 539376 176604 539382 176616
rect 542998 176604 543004 176616
rect 543056 176604 543062 176656
rect 211706 176576 211712 176588
rect 190426 176548 211712 176576
rect 211706 176536 211712 176548
rect 211764 176536 211770 176588
rect 222010 176536 222016 176588
rect 222068 176576 222074 176588
rect 232498 176576 232504 176588
rect 222068 176548 232504 176576
rect 222068 176536 222074 176548
rect 232498 176536 232504 176548
rect 232556 176536 232562 176588
rect 249702 176536 249708 176588
rect 249760 176576 249766 176588
rect 260098 176576 260104 176588
rect 249760 176548 260104 176576
rect 249760 176536 249766 176548
rect 260098 176536 260104 176548
rect 260156 176536 260162 176588
rect 261478 176536 261484 176588
rect 261536 176576 261542 176588
rect 567194 176576 567200 176588
rect 261536 176548 567200 176576
rect 261536 176536 261542 176548
rect 567194 176536 567200 176548
rect 567252 176536 567258 176588
rect 25682 176468 25688 176520
rect 25740 176508 25746 176520
rect 36998 176508 37004 176520
rect 25740 176480 37004 176508
rect 25740 176468 25746 176480
rect 36998 176468 37004 176480
rect 37056 176468 37062 176520
rect 53650 176468 53656 176520
rect 53708 176508 53714 176520
rect 69658 176508 69664 176520
rect 53708 176480 69664 176508
rect 53708 176468 53714 176480
rect 69658 176468 69664 176480
rect 69716 176468 69722 176520
rect 81986 176468 81992 176520
rect 82044 176508 82050 176520
rect 94498 176508 94504 176520
rect 82044 176480 94504 176508
rect 82044 176468 82050 176480
rect 94498 176468 94504 176480
rect 94556 176468 94562 176520
rect 109678 176468 109684 176520
rect 109736 176508 109742 176520
rect 120718 176508 120724 176520
rect 109736 176480 120724 176508
rect 109736 176468 109742 176480
rect 120718 176468 120724 176480
rect 120776 176468 120782 176520
rect 137646 176468 137652 176520
rect 137704 176508 137710 176520
rect 148318 176508 148324 176520
rect 137704 176480 148324 176508
rect 137704 176468 137710 176480
rect 148318 176468 148324 176480
rect 148376 176468 148382 176520
rect 193674 176468 193680 176520
rect 193732 176508 193738 176520
rect 204898 176508 204904 176520
rect 193732 176480 204904 176508
rect 193732 176468 193738 176480
rect 204898 176468 204904 176480
rect 204956 176468 204962 176520
rect 238846 176468 238852 176520
rect 238904 176508 238910 176520
rect 268010 176508 268016 176520
rect 238904 176480 268016 176508
rect 238904 176468 238910 176480
rect 268010 176468 268016 176480
rect 268068 176468 268074 176520
rect 277670 176468 277676 176520
rect 277728 176508 277734 176520
rect 289078 176508 289084 176520
rect 277728 176480 289084 176508
rect 277728 176468 277734 176480
rect 289078 176468 289084 176480
rect 289136 176468 289142 176520
rect 306006 176468 306012 176520
rect 306064 176508 306070 176520
rect 316678 176508 316684 176520
rect 306064 176480 316684 176508
rect 306064 176468 306070 176480
rect 316678 176468 316684 176480
rect 316736 176468 316742 176520
rect 323026 176468 323032 176520
rect 323084 176508 323090 176520
rect 352006 176508 352012 176520
rect 323084 176480 352012 176508
rect 323084 176468 323090 176480
rect 352006 176468 352012 176480
rect 352064 176468 352070 176520
rect 361666 176468 361672 176520
rect 361724 176508 361730 176520
rect 373258 176508 373264 176520
rect 361724 176480 373264 176508
rect 361724 176468 361730 176480
rect 373258 176468 373264 176480
rect 373316 176468 373322 176520
rect 379606 176468 379612 176520
rect 379664 176508 379670 176520
rect 408034 176508 408040 176520
rect 379664 176480 408040 176508
rect 379664 176468 379670 176480
rect 408034 176468 408040 176480
rect 408092 176468 408098 176520
rect 417694 176468 417700 176520
rect 417752 176508 417758 176520
rect 428550 176508 428556 176520
rect 417752 176480 428556 176508
rect 417752 176468 417758 176480
rect 428550 176468 428556 176480
rect 428608 176468 428614 176520
rect 434806 176468 434812 176520
rect 434864 176508 434870 176520
rect 463694 176508 463700 176520
rect 434864 176480 463700 176508
rect 434864 176468 434870 176480
rect 463694 176468 463700 176480
rect 463752 176468 463758 176520
rect 473998 176468 474004 176520
rect 474056 176508 474062 176520
rect 485038 176508 485044 176520
rect 474056 176480 485044 176508
rect 474056 176468 474062 176480
rect 485038 176468 485044 176480
rect 485096 176468 485102 176520
rect 501690 176468 501696 176520
rect 501748 176508 501754 176520
rect 512638 176508 512644 176520
rect 501748 176480 512644 176508
rect 501748 176468 501754 176480
rect 512638 176468 512644 176480
rect 512696 176468 512702 176520
rect 518986 176468 518992 176520
rect 519044 176508 519050 176520
rect 547874 176508 547880 176520
rect 519044 176480 547880 176508
rect 519044 176468 519050 176480
rect 547874 176468 547880 176480
rect 547932 176468 547938 176520
rect 333698 176400 333704 176452
rect 333756 176440 333762 176452
rect 344278 176440 344284 176452
rect 333756 176412 344284 176440
rect 333756 176400 333762 176412
rect 344278 176400 344284 176412
rect 344336 176400 344342 176452
rect 390002 176400 390008 176452
rect 390060 176440 390066 176452
rect 400858 176440 400864 176452
rect 390060 176412 400864 176440
rect 390060 176400 390066 176412
rect 400858 176400 400864 176412
rect 400916 176400 400922 176452
rect 445662 176400 445668 176452
rect 445720 176440 445726 176452
rect 456058 176440 456064 176452
rect 445720 176412 456064 176440
rect 445720 176400 445726 176412
rect 456058 176400 456064 176412
rect 456116 176400 456122 176452
rect 529658 176400 529664 176452
rect 529716 176440 529722 176452
rect 540238 176440 540244 176452
rect 529716 176412 540244 176440
rect 529716 176400 529722 176412
rect 540238 176400 540244 176412
rect 540296 176400 540302 176452
rect 36814 176332 36820 176384
rect 36872 176372 36878 176384
rect 557534 176372 557540 176384
rect 36872 176344 557540 176372
rect 36872 176332 36878 176344
rect 557534 176332 557540 176344
rect 557592 176332 557598 176384
rect 16022 173136 16028 173188
rect 16080 173176 16086 173188
rect 547874 173176 547880 173188
rect 16080 173148 547880 173176
rect 16080 173136 16086 173148
rect 547874 173136 547880 173148
rect 547932 173136 547938 173188
rect 212258 172728 212264 172780
rect 212316 172768 212322 172780
rect 232682 172768 232688 172780
rect 212316 172740 232688 172768
rect 212316 172728 212322 172740
rect 232682 172728 232688 172740
rect 232740 172728 232746 172780
rect 296346 172728 296352 172780
rect 296404 172768 296410 172780
rect 316770 172768 316776 172780
rect 296404 172740 316776 172768
rect 296404 172728 296410 172740
rect 316770 172728 316776 172740
rect 316828 172728 316834 172780
rect 408034 172728 408040 172780
rect 408092 172768 408098 172780
rect 428642 172768 428648 172780
rect 408092 172740 428648 172768
rect 408092 172728 408098 172740
rect 428642 172728 428648 172740
rect 428700 172728 428706 172780
rect 492030 172728 492036 172780
rect 492088 172768 492094 172780
rect 512730 172768 512736 172780
rect 492088 172740 512736 172768
rect 492088 172728 492094 172740
rect 512730 172728 512736 172740
rect 512788 172728 512794 172780
rect 25682 172660 25688 172712
rect 25740 172700 25746 172712
rect 39298 172700 39304 172712
rect 25740 172672 39304 172700
rect 25740 172660 25746 172672
rect 39298 172660 39304 172672
rect 39356 172660 39362 172712
rect 148410 172660 148416 172712
rect 148468 172700 148474 172712
rect 165614 172700 165620 172712
rect 148468 172672 165620 172700
rect 148468 172660 148474 172672
rect 165614 172660 165620 172672
rect 165672 172660 165678 172712
rect 175458 172660 175464 172712
rect 175516 172700 175522 172712
rect 193674 172700 193680 172712
rect 175516 172672 193680 172700
rect 175516 172660 175522 172672
rect 193674 172660 193680 172672
rect 193732 172660 193738 172712
rect 203518 172660 203524 172712
rect 203576 172700 203582 172712
rect 221366 172700 221372 172712
rect 203576 172672 221372 172700
rect 203576 172660 203582 172672
rect 221366 172660 221372 172672
rect 221424 172660 221430 172712
rect 260190 172660 260196 172712
rect 260248 172700 260254 172712
rect 277670 172700 277676 172712
rect 260248 172672 277676 172700
rect 260248 172660 260254 172672
rect 277670 172660 277676 172672
rect 277728 172660 277734 172712
rect 287514 172660 287520 172712
rect 287572 172700 287578 172712
rect 305362 172700 305368 172712
rect 287572 172672 305368 172700
rect 287572 172660 287578 172672
rect 305362 172660 305368 172672
rect 305420 172660 305426 172712
rect 345658 172660 345664 172712
rect 345716 172700 345722 172712
rect 361666 172700 361672 172712
rect 345716 172672 361672 172700
rect 345716 172660 345722 172672
rect 361666 172660 361672 172672
rect 361724 172660 361730 172712
rect 371510 172660 371516 172712
rect 371568 172700 371574 172712
rect 389358 172700 389364 172712
rect 371568 172672 389364 172700
rect 371568 172660 371574 172672
rect 389358 172660 389364 172672
rect 389416 172660 389422 172712
rect 399478 172660 399484 172712
rect 399536 172700 399542 172712
rect 417694 172700 417700 172712
rect 399536 172672 417700 172700
rect 399536 172660 399542 172672
rect 417694 172660 417700 172672
rect 417752 172660 417758 172712
rect 456150 172660 456156 172712
rect 456208 172700 456214 172712
rect 473538 172700 473544 172712
rect 456208 172672 473544 172700
rect 456208 172660 456214 172672
rect 473538 172660 473544 172672
rect 473596 172660 473602 172712
rect 483474 172660 483480 172712
rect 483532 172700 483538 172712
rect 501690 172700 501696 172712
rect 483532 172672 501696 172700
rect 483532 172660 483538 172672
rect 501690 172660 501696 172672
rect 501748 172660 501754 172712
rect 36998 172592 37004 172644
rect 37056 172632 37062 172644
rect 53650 172632 53656 172644
rect 37056 172604 53656 172632
rect 37056 172592 37062 172604
rect 53650 172592 53656 172604
rect 53708 172592 53714 172644
rect 64322 172592 64328 172644
rect 64380 172632 64386 172644
rect 81434 172632 81440 172644
rect 64380 172604 81440 172632
rect 64380 172592 64386 172604
rect 81434 172592 81440 172604
rect 81492 172592 81498 172644
rect 91462 172592 91468 172644
rect 91520 172632 91526 172644
rect 109678 172632 109684 172644
rect 91520 172604 109684 172632
rect 91520 172592 91526 172604
rect 109678 172592 109684 172604
rect 109736 172592 109742 172644
rect 119430 172592 119436 172644
rect 119488 172632 119494 172644
rect 137646 172632 137652 172644
rect 119488 172604 137652 172632
rect 119488 172592 119494 172604
rect 137646 172592 137652 172604
rect 137704 172592 137710 172644
rect 156322 172592 156328 172644
rect 156380 172632 156386 172644
rect 178678 172632 178684 172644
rect 156380 172604 178684 172632
rect 156380 172592 156386 172604
rect 178678 172592 178684 172604
rect 178736 172592 178742 172644
rect 232590 172592 232596 172644
rect 232648 172632 232654 172644
rect 249702 172632 249708 172644
rect 232648 172604 249708 172632
rect 232648 172592 232654 172604
rect 249702 172592 249708 172604
rect 249760 172592 249766 172644
rect 268010 172592 268016 172644
rect 268068 172632 268074 172644
rect 287698 172632 287704 172644
rect 268068 172604 287704 172632
rect 268068 172592 268074 172604
rect 287698 172592 287704 172604
rect 287756 172592 287762 172644
rect 315482 172592 315488 172644
rect 315540 172632 315546 172644
rect 333698 172632 333704 172644
rect 315540 172604 333704 172632
rect 315540 172592 315546 172604
rect 333698 172592 333704 172604
rect 333756 172592 333762 172644
rect 352006 172592 352012 172644
rect 352064 172632 352070 172644
rect 374638 172632 374644 172644
rect 352064 172604 374644 172632
rect 352064 172592 352070 172604
rect 374638 172592 374644 172604
rect 374696 172592 374702 172644
rect 428458 172592 428464 172644
rect 428516 172632 428522 172644
rect 445662 172632 445668 172644
rect 428516 172604 445668 172632
rect 428516 172592 428522 172604
rect 445662 172592 445668 172604
rect 445720 172592 445726 172644
rect 464338 172592 464344 172644
rect 464396 172632 464402 172644
rect 483658 172632 483664 172644
rect 464396 172604 483664 172632
rect 464396 172592 464402 172604
rect 483658 172592 483664 172604
rect 483716 172592 483722 172644
rect 511442 172592 511448 172644
rect 511500 172632 511506 172644
rect 529658 172632 529664 172644
rect 511500 172604 529664 172632
rect 511500 172592 511506 172604
rect 529658 172592 529664 172604
rect 529716 172592 529722 172644
rect 542998 172592 543004 172644
rect 543056 172632 543062 172644
rect 557534 172632 557540 172644
rect 543056 172604 557540 172632
rect 543056 172592 543062 172604
rect 557534 172592 557540 172604
rect 557592 172592 557598 172644
rect 36906 172524 36912 172576
rect 36964 172564 36970 172576
rect 63310 172564 63316 172576
rect 36964 172536 63316 172564
rect 36964 172524 36970 172536
rect 63310 172524 63316 172536
rect 63368 172524 63374 172576
rect 66898 172524 66904 172576
rect 66956 172564 66962 172576
rect 91094 172564 91100 172576
rect 66956 172536 91100 172564
rect 66956 172524 66962 172536
rect 91094 172524 91100 172536
rect 91152 172524 91158 172576
rect 94498 172524 94504 172576
rect 94556 172564 94562 172576
rect 119338 172564 119344 172576
rect 94556 172536 119344 172564
rect 94556 172524 94562 172536
rect 119338 172524 119344 172536
rect 119396 172524 119402 172576
rect 120718 172524 120724 172576
rect 120776 172564 120782 172576
rect 147306 172564 147312 172576
rect 120776 172536 147312 172564
rect 120776 172524 120782 172536
rect 147306 172524 147312 172536
rect 147364 172524 147370 172576
rect 148318 172524 148324 172576
rect 148376 172564 148382 172576
rect 175274 172564 175280 172576
rect 148376 172536 175280 172564
rect 148376 172524 148382 172536
rect 175274 172524 175280 172536
rect 175332 172524 175338 172576
rect 177298 172524 177304 172576
rect 177356 172564 177362 172576
rect 203334 172564 203340 172576
rect 177356 172536 203340 172564
rect 177356 172524 177362 172536
rect 203334 172524 203340 172536
rect 203392 172524 203398 172576
rect 204898 172524 204904 172576
rect 204956 172564 204962 172576
rect 231026 172564 231032 172576
rect 204956 172536 231032 172564
rect 204956 172524 204962 172536
rect 231026 172524 231032 172536
rect 231084 172524 231090 172576
rect 232498 172524 232504 172576
rect 232556 172564 232562 172576
rect 259362 172564 259368 172576
rect 232556 172536 259368 172564
rect 232556 172524 232562 172536
rect 259362 172524 259368 172536
rect 259420 172524 259426 172576
rect 260098 172524 260104 172576
rect 260156 172564 260162 172576
rect 287330 172564 287336 172576
rect 260156 172536 287336 172564
rect 260156 172524 260162 172536
rect 287330 172524 287336 172536
rect 287388 172524 287394 172576
rect 289078 172524 289084 172576
rect 289136 172564 289142 172576
rect 315022 172564 315028 172576
rect 289136 172536 315028 172564
rect 289136 172524 289142 172536
rect 315022 172524 315028 172536
rect 315080 172524 315086 172576
rect 316678 172524 316684 172576
rect 316736 172564 316742 172576
rect 343358 172564 343364 172576
rect 316736 172536 343364 172564
rect 316736 172524 316742 172536
rect 343358 172524 343364 172536
rect 343416 172524 343422 172576
rect 344278 172524 344284 172576
rect 344336 172564 344342 172576
rect 371326 172564 371332 172576
rect 344336 172536 371332 172564
rect 344336 172524 344342 172536
rect 371326 172524 371332 172536
rect 371384 172524 371390 172576
rect 373258 172524 373264 172576
rect 373316 172564 373322 172576
rect 399018 172564 399024 172576
rect 373316 172536 399024 172564
rect 373316 172524 373322 172536
rect 399018 172524 399024 172536
rect 399076 172524 399082 172576
rect 400858 172524 400864 172576
rect 400916 172564 400922 172576
rect 427354 172564 427360 172576
rect 400916 172536 427360 172564
rect 400916 172524 400922 172536
rect 427354 172524 427360 172536
rect 427412 172524 427418 172576
rect 428550 172524 428556 172576
rect 428608 172564 428614 172576
rect 455322 172564 455328 172576
rect 428608 172536 455328 172564
rect 428608 172524 428614 172536
rect 455322 172524 455328 172536
rect 455380 172524 455386 172576
rect 456058 172524 456064 172576
rect 456116 172564 456122 172576
rect 483198 172564 483204 172576
rect 456116 172536 483204 172564
rect 456116 172524 456122 172536
rect 483198 172524 483204 172536
rect 483256 172524 483262 172576
rect 485038 172524 485044 172576
rect 485096 172564 485102 172576
rect 511350 172564 511356 172576
rect 485096 172536 511356 172564
rect 485096 172524 485102 172536
rect 511350 172524 511356 172536
rect 511408 172524 511414 172576
rect 512638 172524 512644 172576
rect 512696 172564 512702 172576
rect 539318 172564 539324 172576
rect 512696 172536 539324 172564
rect 512696 172524 512702 172536
rect 539318 172524 539324 172536
rect 539376 172524 539382 172576
rect 540238 172524 540244 172576
rect 540296 172564 540302 172576
rect 567194 172564 567200 172576
rect 540296 172536 567200 172564
rect 540296 172524 540302 172536
rect 567194 172524 567200 172536
rect 567252 172524 567258 172576
rect 37918 170348 37924 170400
rect 37976 170388 37982 170400
rect 545758 170388 545764 170400
rect 37976 170360 545764 170388
rect 37976 170348 37982 170360
rect 545758 170348 545764 170360
rect 545816 170348 545822 170400
rect 35618 169736 35624 169788
rect 35676 169776 35682 169788
rect 36814 169776 36820 169788
rect 35676 169748 36820 169776
rect 35676 169736 35682 169748
rect 36814 169736 36820 169748
rect 36872 169736 36878 169788
rect 63586 156612 63592 156664
rect 63644 156652 63650 156664
rect 64322 156652 64328 156664
rect 63644 156624 64328 156652
rect 63644 156612 63650 156624
rect 64322 156612 64328 156624
rect 64380 156612 64386 156664
rect 147674 156612 147680 156664
rect 147732 156652 147738 156664
rect 148410 156652 148416 156664
rect 147732 156624 148416 156652
rect 147732 156612 147738 156624
rect 148410 156612 148416 156624
rect 148468 156612 148474 156664
rect 259730 156612 259736 156664
rect 259788 156652 259794 156664
rect 260190 156652 260196 156664
rect 259788 156624 260196 156652
rect 259788 156612 259794 156624
rect 260190 156612 260196 156624
rect 260248 156612 260254 156664
rect 455690 156612 455696 156664
rect 455748 156652 455754 156664
rect 456150 156652 456156 156664
rect 455748 156624 456156 156652
rect 455748 156612 455754 156624
rect 456150 156612 456156 156624
rect 456208 156612 456214 156664
rect 287698 153144 287704 153196
rect 287756 153184 287762 153196
rect 295702 153184 295708 153196
rect 287756 153156 295708 153184
rect 287756 153144 287762 153156
rect 295702 153144 295708 153156
rect 295760 153144 295766 153196
rect 316770 153144 316776 153196
rect 316828 153184 316834 153196
rect 323670 153184 323676 153196
rect 316828 153156 323676 153184
rect 316828 153144 316834 153156
rect 323670 153144 323676 153156
rect 323728 153144 323734 153196
rect 232682 152532 232688 152584
rect 232740 152572 232746 152584
rect 239766 152572 239772 152584
rect 232740 152544 239772 152572
rect 232740 152532 232746 152544
rect 239766 152532 239772 152544
rect 239824 152532 239830 152584
rect 428642 152464 428648 152516
rect 428700 152504 428706 152516
rect 435726 152504 435732 152516
rect 428700 152476 435732 152504
rect 428700 152464 428706 152476
rect 435726 152464 435732 152476
rect 435784 152464 435790 152516
rect 483658 152464 483664 152516
rect 483716 152504 483722 152516
rect 491662 152504 491668 152516
rect 483716 152476 491668 152504
rect 483716 152464 483722 152476
rect 491662 152464 491668 152476
rect 491720 152464 491726 152516
rect 512730 152192 512736 152244
rect 512788 152232 512794 152244
rect 519630 152232 519636 152244
rect 512788 152204 519636 152232
rect 512788 152192 512794 152204
rect 519630 152192 519636 152204
rect 519688 152192 519694 152244
rect 13722 151716 13728 151768
rect 13780 151756 13786 151768
rect 66254 151756 66260 151768
rect 13780 151728 66260 151756
rect 13780 151716 13786 151728
rect 66254 151716 66260 151728
rect 66312 151716 66318 151768
rect 70302 151716 70308 151768
rect 70360 151756 70366 151768
rect 121454 151756 121460 151768
rect 70360 151728 121460 151756
rect 70360 151716 70366 151728
rect 121454 151716 121460 151728
rect 121512 151716 121518 151768
rect 126882 151716 126888 151768
rect 126940 151756 126946 151768
rect 178034 151756 178040 151768
rect 126940 151728 178040 151756
rect 126940 151716 126946 151728
rect 178034 151716 178040 151728
rect 178092 151716 178098 151768
rect 209682 151716 209688 151768
rect 209740 151756 209746 151768
rect 262214 151756 262220 151768
rect 209740 151728 262220 151756
rect 209740 151716 209746 151728
rect 262214 151716 262220 151728
rect 262272 151716 262278 151768
rect 266262 151716 266268 151768
rect 266320 151756 266326 151768
rect 317414 151756 317420 151768
rect 266320 151728 317420 151756
rect 266320 151716 266326 151728
rect 317414 151716 317420 151728
rect 317472 151716 317478 151768
rect 322842 151716 322848 151768
rect 322900 151756 322906 151768
rect 373994 151756 374000 151768
rect 322900 151728 374000 151756
rect 322900 151716 322906 151728
rect 373994 151716 374000 151728
rect 374052 151716 374058 151768
rect 405642 151716 405648 151768
rect 405700 151756 405706 151768
rect 458174 151756 458180 151768
rect 405700 151728 458180 151756
rect 405700 151716 405706 151728
rect 458174 151716 458180 151728
rect 458232 151716 458238 151768
rect 489822 151716 489828 151768
rect 489880 151756 489886 151768
rect 542354 151756 542360 151768
rect 489880 151728 542360 151756
rect 489880 151716 489886 151728
rect 542354 151716 542360 151728
rect 542412 151716 542418 151768
rect 35618 151648 35624 151700
rect 35676 151688 35682 151700
rect 36998 151688 37004 151700
rect 35676 151660 37004 151688
rect 35676 151648 35682 151660
rect 36998 151648 37004 151660
rect 37056 151648 37062 151700
rect 42702 151648 42708 151700
rect 42760 151688 42766 151700
rect 93854 151688 93860 151700
rect 42760 151660 93860 151688
rect 42760 151648 42766 151660
rect 93854 151648 93860 151660
rect 93912 151648 93918 151700
rect 97902 151648 97908 151700
rect 97960 151688 97966 151700
rect 149054 151688 149060 151700
rect 97960 151660 149060 151688
rect 97960 151648 97966 151660
rect 149054 151648 149060 151660
rect 149112 151648 149118 151700
rect 154482 151648 154488 151700
rect 154540 151688 154546 151700
rect 205634 151688 205640 151700
rect 154540 151660 205640 151688
rect 154540 151648 154546 151660
rect 205634 151648 205640 151660
rect 205692 151648 205698 151700
rect 231670 151648 231676 151700
rect 231728 151688 231734 151700
rect 232590 151688 232596 151700
rect 231728 151660 232596 151688
rect 231728 151648 231734 151660
rect 232590 151648 232596 151660
rect 232648 151648 232654 151700
rect 238662 151648 238668 151700
rect 238720 151688 238726 151700
rect 289814 151688 289820 151700
rect 238720 151660 289820 151688
rect 238720 151648 238726 151660
rect 289814 151648 289820 151660
rect 289872 151648 289878 151700
rect 293862 151648 293868 151700
rect 293920 151688 293926 151700
rect 293920 151660 335354 151688
rect 293920 151648 293926 151660
rect 182082 151580 182088 151632
rect 182140 151620 182146 151632
rect 233234 151620 233240 151632
rect 182140 151592 233240 151620
rect 182140 151580 182146 151592
rect 233234 151580 233240 151592
rect 233292 151580 233298 151632
rect 335326 151620 335354 151660
rect 343634 151648 343640 151700
rect 343692 151688 343698 151700
rect 345658 151688 345664 151700
rect 343692 151660 345664 151688
rect 343692 151648 343698 151660
rect 345658 151648 345664 151660
rect 345716 151648 345722 151700
rect 350442 151648 350448 151700
rect 350500 151688 350506 151700
rect 401594 151688 401600 151700
rect 350500 151660 401600 151688
rect 350500 151648 350506 151660
rect 401594 151648 401600 151660
rect 401652 151648 401658 151700
rect 434622 151648 434628 151700
rect 434680 151688 434686 151700
rect 485774 151688 485780 151700
rect 434680 151660 485780 151688
rect 434680 151648 434686 151660
rect 485774 151648 485780 151660
rect 485832 151648 485838 151700
rect 518802 151648 518808 151700
rect 518860 151688 518866 151700
rect 569954 151688 569960 151700
rect 518860 151660 569960 151688
rect 518860 151648 518866 151660
rect 569954 151648 569960 151660
rect 570012 151648 570018 151700
rect 345014 151620 345020 151632
rect 335326 151592 345020 151620
rect 345014 151580 345020 151592
rect 345072 151580 345078 151632
rect 378042 151580 378048 151632
rect 378100 151620 378106 151632
rect 429194 151620 429200 151632
rect 378100 151592 429200 151620
rect 378100 151580 378106 151592
rect 429194 151580 429200 151592
rect 429252 151580 429258 151632
rect 462222 151580 462228 151632
rect 462280 151620 462286 151632
rect 513374 151620 513380 151632
rect 462280 151592 513380 151620
rect 462280 151580 462286 151592
rect 513374 151580 513380 151592
rect 513432 151580 513438 151632
rect 539502 151580 539508 151632
rect 539560 151620 539566 151632
rect 542998 151620 543004 151632
rect 539560 151592 543004 151620
rect 539560 151580 539566 151592
rect 542998 151580 543004 151592
rect 543056 151580 543062 151632
rect 178678 148996 178684 149048
rect 178736 149036 178742 149048
rect 184014 149036 184020 149048
rect 178736 149008 184020 149036
rect 178736 148996 178742 149008
rect 184014 148996 184020 149008
rect 184072 148996 184078 149048
rect 374638 148996 374644 149048
rect 374696 149036 374702 149048
rect 379698 149036 379704 149048
rect 374696 149008 379704 149036
rect 374696 148996 374702 149008
rect 379698 148996 379704 149008
rect 379756 148996 379762 149048
rect 15194 148928 15200 148980
rect 15252 148968 15258 148980
rect 43990 148968 43996 148980
rect 15252 148940 43996 148968
rect 15252 148928 15258 148940
rect 43990 148928 43996 148940
rect 44048 148928 44054 148980
rect 71038 148928 71044 148980
rect 71096 148968 71102 148980
rect 567194 148968 567200 148980
rect 71096 148940 567200 148968
rect 71096 148928 71102 148940
rect 567194 148928 567200 148940
rect 567252 148928 567258 148980
rect 25682 148860 25688 148912
rect 25740 148900 25746 148912
rect 36906 148900 36912 148912
rect 25740 148872 36912 148900
rect 25740 148860 25746 148872
rect 36906 148860 36912 148872
rect 36964 148860 36970 148912
rect 53650 148860 53656 148912
rect 53708 148900 53714 148912
rect 66898 148900 66904 148912
rect 53708 148872 66904 148900
rect 53708 148860 53714 148872
rect 66898 148860 66904 148872
rect 66956 148860 66962 148912
rect 71866 148860 71872 148912
rect 71924 148900 71930 148912
rect 100018 148900 100024 148912
rect 71924 148872 100024 148900
rect 71924 148860 71930 148872
rect 100018 148860 100024 148872
rect 100076 148860 100082 148912
rect 127986 148900 127992 148912
rect 103486 148872 127992 148900
rect 42886 148792 42892 148844
rect 42944 148832 42950 148844
rect 72050 148832 72056 148844
rect 42944 148804 72056 148832
rect 42944 148792 42950 148804
rect 72050 148792 72056 148804
rect 72108 148792 72114 148844
rect 81986 148792 81992 148844
rect 82044 148832 82050 148844
rect 94498 148832 94504 148844
rect 82044 148804 94504 148832
rect 82044 148792 82050 148804
rect 94498 148792 94504 148804
rect 94556 148792 94562 148844
rect 99466 148792 99472 148844
rect 99524 148832 99530 148844
rect 103486 148832 103514 148872
rect 127986 148860 127992 148872
rect 128044 148860 128050 148912
rect 156046 148900 156052 148912
rect 132466 148872 156052 148900
rect 99524 148804 103514 148832
rect 99524 148792 99530 148804
rect 109678 148792 109684 148844
rect 109736 148832 109742 148844
rect 120718 148832 120724 148844
rect 109736 148804 120724 148832
rect 109736 148792 109742 148804
rect 120718 148792 120724 148804
rect 120776 148792 120782 148844
rect 127066 148792 127072 148844
rect 127124 148832 127130 148844
rect 132466 148832 132494 148872
rect 156046 148860 156052 148872
rect 156104 148860 156110 148912
rect 165982 148860 165988 148912
rect 166040 148900 166046 148912
rect 177298 148900 177304 148912
rect 166040 148872 177304 148900
rect 166040 148860 166046 148872
rect 177298 148860 177304 148872
rect 177356 148860 177362 148912
rect 183646 148860 183652 148912
rect 183704 148900 183710 148912
rect 211706 148900 211712 148912
rect 183704 148872 211712 148900
rect 183704 148860 183710 148872
rect 211706 148860 211712 148872
rect 211764 148860 211770 148912
rect 222010 148860 222016 148912
rect 222068 148900 222074 148912
rect 232498 148900 232504 148912
rect 222068 148872 232504 148900
rect 222068 148860 222074 148872
rect 232498 148860 232504 148872
rect 232556 148860 232562 148912
rect 238846 148860 238852 148912
rect 238904 148900 238910 148912
rect 268010 148900 268016 148912
rect 238904 148872 268016 148900
rect 238904 148860 238910 148872
rect 268010 148860 268016 148872
rect 268068 148860 268074 148912
rect 277670 148860 277676 148912
rect 277728 148900 277734 148912
rect 289078 148900 289084 148912
rect 277728 148872 289084 148900
rect 277728 148860 277734 148872
rect 289078 148860 289084 148872
rect 289136 148860 289142 148912
rect 306006 148860 306012 148912
rect 306064 148900 306070 148912
rect 316678 148900 316684 148912
rect 306064 148872 316684 148900
rect 306064 148860 306070 148872
rect 316678 148860 316684 148872
rect 316736 148860 316742 148912
rect 323026 148860 323032 148912
rect 323084 148900 323090 148912
rect 352006 148900 352012 148912
rect 323084 148872 352012 148900
rect 323084 148860 323090 148872
rect 352006 148860 352012 148872
rect 352064 148860 352070 148912
rect 361666 148860 361672 148912
rect 361724 148900 361730 148912
rect 373258 148900 373264 148912
rect 361724 148872 373264 148900
rect 361724 148860 361730 148872
rect 373258 148860 373264 148872
rect 373316 148860 373322 148912
rect 379606 148860 379612 148912
rect 379664 148900 379670 148912
rect 408034 148900 408040 148912
rect 379664 148872 408040 148900
rect 379664 148860 379670 148872
rect 408034 148860 408040 148872
rect 408092 148860 408098 148912
rect 417694 148860 417700 148912
rect 417752 148900 417758 148912
rect 428550 148900 428556 148912
rect 417752 148872 428556 148900
rect 417752 148860 417758 148872
rect 428550 148860 428556 148872
rect 428608 148860 428614 148912
rect 434806 148860 434812 148912
rect 434864 148900 434870 148912
rect 463694 148900 463700 148912
rect 434864 148872 463700 148900
rect 434864 148860 434870 148872
rect 463694 148860 463700 148872
rect 463752 148860 463758 148912
rect 473998 148860 474004 148912
rect 474056 148900 474062 148912
rect 485038 148900 485044 148912
rect 474056 148872 485044 148900
rect 474056 148860 474062 148872
rect 485038 148860 485044 148872
rect 485096 148860 485102 148912
rect 501690 148860 501696 148912
rect 501748 148900 501754 148912
rect 512638 148900 512644 148912
rect 501748 148872 512644 148900
rect 501748 148860 501754 148872
rect 512638 148860 512644 148872
rect 512696 148860 512702 148912
rect 518986 148860 518992 148912
rect 519044 148900 519050 148912
rect 547874 148900 547880 148912
rect 519044 148872 547880 148900
rect 519044 148860 519050 148872
rect 547874 148860 547880 148872
rect 547932 148860 547938 148912
rect 127124 148804 132494 148832
rect 127124 148792 127130 148804
rect 137646 148792 137652 148844
rect 137704 148832 137710 148844
rect 148318 148832 148324 148844
rect 137704 148804 148324 148832
rect 137704 148792 137710 148804
rect 148318 148792 148324 148804
rect 148376 148792 148382 148844
rect 193674 148792 193680 148844
rect 193732 148832 193738 148844
rect 204898 148832 204904 148844
rect 193732 148804 204904 148832
rect 193732 148792 193738 148804
rect 204898 148792 204904 148804
rect 204956 148792 204962 148844
rect 249702 148792 249708 148844
rect 249760 148832 249766 148844
rect 260098 148832 260104 148844
rect 249760 148804 260104 148832
rect 249760 148792 249766 148804
rect 260098 148792 260104 148804
rect 260156 148792 260162 148844
rect 333698 148792 333704 148844
rect 333756 148832 333762 148844
rect 344278 148832 344284 148844
rect 333756 148804 344284 148832
rect 333756 148792 333762 148804
rect 344278 148792 344284 148804
rect 344336 148792 344342 148844
rect 390002 148792 390008 148844
rect 390060 148832 390066 148844
rect 400858 148832 400864 148844
rect 390060 148804 400864 148832
rect 390060 148792 390066 148804
rect 400858 148792 400864 148804
rect 400916 148792 400922 148844
rect 445662 148792 445668 148844
rect 445720 148832 445726 148844
rect 456058 148832 456064 148844
rect 445720 148804 456064 148832
rect 445720 148792 445726 148804
rect 456058 148792 456064 148804
rect 456116 148792 456122 148844
rect 529658 148792 529664 148844
rect 529716 148832 529722 148844
rect 540238 148832 540244 148844
rect 529716 148804 540244 148832
rect 529716 148792 529722 148804
rect 540238 148792 540244 148804
rect 540296 148792 540302 148844
rect 36722 148724 36728 148776
rect 36780 148764 36786 148776
rect 557534 148764 557540 148776
rect 36780 148736 557540 148764
rect 36780 148724 36786 148736
rect 557534 148724 557540 148736
rect 557592 148724 557598 148776
rect 16022 146888 16028 146940
rect 16080 146928 16086 146940
rect 547874 146928 547880 146940
rect 16080 146900 547880 146928
rect 16080 146888 16086 146900
rect 547874 146888 547880 146900
rect 547932 146888 547938 146940
rect 25682 146480 25688 146532
rect 25740 146520 25746 146532
rect 71038 146520 71044 146532
rect 25740 146492 71044 146520
rect 25740 146480 25746 146492
rect 71038 146480 71044 146492
rect 71096 146480 71102 146532
rect 212350 146480 212356 146532
rect 212408 146520 212414 146532
rect 232682 146520 232688 146532
rect 212408 146492 232688 146520
rect 212408 146480 212414 146492
rect 232682 146480 232688 146492
rect 232740 146480 232746 146532
rect 296346 146480 296352 146532
rect 296404 146520 296410 146532
rect 316770 146520 316776 146532
rect 296404 146492 316776 146520
rect 296404 146480 296410 146492
rect 316770 146480 316776 146492
rect 316828 146480 316834 146532
rect 408034 146480 408040 146532
rect 408092 146520 408098 146532
rect 428642 146520 428648 146532
rect 408092 146492 428648 146520
rect 408092 146480 408098 146492
rect 428642 146480 428648 146492
rect 428700 146480 428706 146532
rect 492030 146480 492036 146532
rect 492088 146520 492094 146532
rect 512730 146520 512736 146532
rect 492088 146492 512736 146520
rect 492088 146480 492094 146492
rect 512730 146480 512736 146492
rect 512788 146480 512794 146532
rect 36906 146412 36912 146464
rect 36964 146452 36970 146464
rect 53650 146452 53656 146464
rect 36964 146424 53656 146452
rect 36964 146412 36970 146424
rect 53650 146412 53656 146424
rect 53708 146412 53714 146464
rect 148410 146412 148416 146464
rect 148468 146452 148474 146464
rect 165706 146452 165712 146464
rect 148468 146424 165712 146452
rect 148468 146412 148474 146424
rect 165706 146412 165712 146424
rect 165764 146412 165770 146464
rect 175458 146412 175464 146464
rect 175516 146452 175522 146464
rect 193674 146452 193680 146464
rect 175516 146424 193680 146452
rect 175516 146412 175522 146424
rect 193674 146412 193680 146424
rect 193732 146412 193738 146464
rect 203518 146412 203524 146464
rect 203576 146452 203582 146464
rect 221366 146452 221372 146464
rect 203576 146424 221372 146452
rect 203576 146412 203582 146424
rect 221366 146412 221372 146424
rect 221424 146412 221430 146464
rect 260098 146412 260104 146464
rect 260156 146452 260162 146464
rect 277670 146452 277676 146464
rect 260156 146424 277676 146452
rect 260156 146412 260162 146424
rect 277670 146412 277676 146424
rect 277728 146412 277734 146464
rect 287514 146412 287520 146464
rect 287572 146452 287578 146464
rect 305362 146452 305368 146464
rect 287572 146424 305368 146452
rect 287572 146412 287578 146424
rect 305362 146412 305368 146424
rect 305420 146412 305426 146464
rect 345658 146412 345664 146464
rect 345716 146452 345722 146464
rect 361666 146452 361672 146464
rect 345716 146424 361672 146452
rect 345716 146412 345722 146424
rect 361666 146412 361672 146424
rect 361724 146412 361730 146464
rect 371510 146412 371516 146464
rect 371568 146452 371574 146464
rect 389358 146452 389364 146464
rect 371568 146424 389364 146452
rect 371568 146412 371574 146424
rect 389358 146412 389364 146424
rect 389416 146412 389422 146464
rect 399478 146412 399484 146464
rect 399536 146452 399542 146464
rect 417694 146452 417700 146464
rect 399536 146424 417700 146452
rect 399536 146412 399542 146424
rect 417694 146412 417700 146424
rect 417752 146412 417758 146464
rect 456058 146412 456064 146464
rect 456116 146452 456122 146464
rect 473354 146452 473360 146464
rect 456116 146424 473360 146452
rect 456116 146412 456122 146424
rect 473354 146412 473360 146424
rect 473412 146412 473418 146464
rect 483474 146412 483480 146464
rect 483532 146452 483538 146464
rect 501690 146452 501696 146464
rect 483532 146424 501696 146452
rect 483532 146412 483538 146424
rect 501690 146412 501696 146424
rect 501748 146412 501754 146464
rect 36998 146344 37004 146396
rect 37056 146384 37062 146396
rect 63310 146384 63316 146396
rect 37056 146356 63316 146384
rect 37056 146344 37062 146356
rect 63310 146344 63316 146356
rect 63368 146344 63374 146396
rect 64322 146344 64328 146396
rect 64380 146384 64386 146396
rect 81434 146384 81440 146396
rect 64380 146356 81440 146384
rect 64380 146344 64386 146356
rect 81434 146344 81440 146356
rect 81492 146344 81498 146396
rect 91462 146344 91468 146396
rect 91520 146384 91526 146396
rect 109678 146384 109684 146396
rect 91520 146356 109684 146384
rect 91520 146344 91526 146356
rect 109678 146344 109684 146356
rect 109736 146344 109742 146396
rect 119430 146344 119436 146396
rect 119488 146384 119494 146396
rect 137646 146384 137652 146396
rect 119488 146356 137652 146384
rect 119488 146344 119494 146356
rect 137646 146344 137652 146356
rect 137704 146344 137710 146396
rect 156322 146344 156328 146396
rect 156380 146384 156386 146396
rect 178678 146384 178684 146396
rect 156380 146356 178684 146384
rect 156380 146344 156386 146356
rect 178678 146344 178684 146356
rect 178736 146344 178742 146396
rect 232498 146344 232504 146396
rect 232556 146384 232562 146396
rect 249702 146384 249708 146396
rect 232556 146356 249708 146384
rect 232556 146344 232562 146356
rect 249702 146344 249708 146356
rect 249760 146344 249766 146396
rect 268010 146344 268016 146396
rect 268068 146384 268074 146396
rect 287698 146384 287704 146396
rect 268068 146356 287704 146384
rect 268068 146344 268074 146356
rect 287698 146344 287704 146356
rect 287756 146344 287762 146396
rect 315482 146344 315488 146396
rect 315540 146384 315546 146396
rect 333698 146384 333704 146396
rect 315540 146356 333704 146384
rect 315540 146344 315546 146356
rect 333698 146344 333704 146356
rect 333756 146344 333762 146396
rect 352006 146344 352012 146396
rect 352064 146384 352070 146396
rect 374638 146384 374644 146396
rect 352064 146356 374644 146384
rect 352064 146344 352070 146356
rect 374638 146344 374644 146356
rect 374696 146344 374702 146396
rect 428458 146344 428464 146396
rect 428516 146384 428522 146396
rect 445662 146384 445668 146396
rect 428516 146356 445668 146384
rect 428516 146344 428522 146356
rect 445662 146344 445668 146356
rect 445720 146344 445726 146396
rect 464338 146344 464344 146396
rect 464396 146384 464402 146396
rect 483658 146384 483664 146396
rect 464396 146356 483664 146384
rect 464396 146344 464402 146356
rect 483658 146344 483664 146356
rect 483716 146344 483722 146396
rect 511442 146344 511448 146396
rect 511500 146384 511506 146396
rect 529658 146384 529664 146396
rect 511500 146356 529664 146384
rect 511500 146344 511506 146356
rect 529658 146344 529664 146356
rect 529716 146344 529722 146396
rect 542998 146344 543004 146396
rect 543056 146384 543062 146396
rect 557534 146384 557540 146396
rect 543056 146356 557540 146384
rect 543056 146344 543062 146356
rect 557534 146344 557540 146356
rect 557592 146344 557598 146396
rect 69658 146276 69664 146328
rect 69716 146316 69722 146328
rect 91094 146316 91100 146328
rect 69716 146288 91100 146316
rect 69716 146276 69722 146288
rect 91094 146276 91100 146288
rect 91152 146276 91158 146328
rect 94498 146276 94504 146328
rect 94556 146316 94562 146328
rect 119338 146316 119344 146328
rect 94556 146288 119344 146316
rect 94556 146276 94562 146288
rect 119338 146276 119344 146288
rect 119396 146276 119402 146328
rect 120718 146276 120724 146328
rect 120776 146316 120782 146328
rect 147306 146316 147312 146328
rect 120776 146288 147312 146316
rect 120776 146276 120782 146288
rect 147306 146276 147312 146288
rect 147364 146276 147370 146328
rect 148318 146276 148324 146328
rect 148376 146316 148382 146328
rect 175366 146316 175372 146328
rect 148376 146288 175372 146316
rect 148376 146276 148382 146288
rect 175366 146276 175372 146288
rect 175424 146276 175430 146328
rect 177298 146276 177304 146328
rect 177356 146316 177362 146328
rect 203334 146316 203340 146328
rect 177356 146288 203340 146316
rect 177356 146276 177362 146288
rect 203334 146276 203340 146288
rect 203392 146276 203398 146328
rect 204898 146276 204904 146328
rect 204956 146316 204962 146328
rect 231026 146316 231032 146328
rect 204956 146288 231032 146316
rect 204956 146276 204962 146288
rect 231026 146276 231032 146288
rect 231084 146276 231090 146328
rect 232590 146276 232596 146328
rect 232648 146316 232654 146328
rect 259362 146316 259368 146328
rect 232648 146288 259368 146316
rect 232648 146276 232654 146288
rect 259362 146276 259368 146288
rect 259420 146276 259426 146328
rect 260190 146276 260196 146328
rect 260248 146316 260254 146328
rect 287330 146316 287336 146328
rect 260248 146288 287336 146316
rect 260248 146276 260254 146288
rect 287330 146276 287336 146288
rect 287388 146276 287394 146328
rect 289078 146276 289084 146328
rect 289136 146316 289142 146328
rect 315022 146316 315028 146328
rect 289136 146288 315028 146316
rect 289136 146276 289142 146288
rect 315022 146276 315028 146288
rect 315080 146276 315086 146328
rect 316678 146276 316684 146328
rect 316736 146316 316742 146328
rect 343358 146316 343364 146328
rect 316736 146288 343364 146316
rect 316736 146276 316742 146288
rect 343358 146276 343364 146288
rect 343416 146276 343422 146328
rect 344278 146276 344284 146328
rect 344336 146316 344342 146328
rect 371326 146316 371332 146328
rect 344336 146288 371332 146316
rect 344336 146276 344342 146288
rect 371326 146276 371332 146288
rect 371384 146276 371390 146328
rect 373258 146276 373264 146328
rect 373316 146316 373322 146328
rect 399018 146316 399024 146328
rect 373316 146288 399024 146316
rect 373316 146276 373322 146288
rect 399018 146276 399024 146288
rect 399076 146276 399082 146328
rect 400858 146276 400864 146328
rect 400916 146316 400922 146328
rect 427354 146316 427360 146328
rect 400916 146288 427360 146316
rect 400916 146276 400922 146288
rect 427354 146276 427360 146288
rect 427412 146276 427418 146328
rect 428550 146276 428556 146328
rect 428608 146316 428614 146328
rect 455322 146316 455328 146328
rect 428608 146288 455328 146316
rect 428608 146276 428614 146288
rect 455322 146276 455328 146288
rect 455380 146276 455386 146328
rect 456150 146276 456156 146328
rect 456208 146316 456214 146328
rect 483014 146316 483020 146328
rect 456208 146288 483020 146316
rect 456208 146276 456214 146288
rect 483014 146276 483020 146288
rect 483072 146276 483078 146328
rect 485038 146276 485044 146328
rect 485096 146316 485102 146328
rect 511350 146316 511356 146328
rect 485096 146288 511356 146316
rect 485096 146276 485102 146288
rect 511350 146276 511356 146288
rect 511408 146276 511414 146328
rect 512638 146276 512644 146328
rect 512696 146316 512702 146328
rect 539318 146316 539324 146328
rect 512696 146288 539324 146316
rect 512696 146276 512702 146288
rect 539318 146276 539324 146288
rect 539376 146276 539382 146328
rect 540238 146276 540244 146328
rect 540296 146316 540302 146328
rect 567194 146316 567200 146328
rect 540296 146288 567200 146316
rect 540296 146276 540302 146288
rect 567194 146276 567200 146288
rect 567252 146276 567258 146328
rect 37918 144168 37924 144220
rect 37976 144208 37982 144220
rect 545758 144208 545764 144220
rect 37976 144180 545764 144208
rect 37976 144168 37982 144180
rect 545758 144168 545764 144180
rect 545816 144168 545822 144220
rect 35618 143556 35624 143608
rect 35676 143596 35682 143608
rect 36722 143596 36728 143608
rect 35676 143568 36728 143596
rect 35676 143556 35682 143568
rect 36722 143556 36728 143568
rect 36780 143556 36786 143608
rect 63586 128256 63592 128308
rect 63644 128296 63650 128308
rect 64322 128296 64328 128308
rect 63644 128268 64328 128296
rect 63644 128256 63650 128268
rect 64322 128256 64328 128268
rect 64380 128256 64386 128308
rect 147674 128256 147680 128308
rect 147732 128296 147738 128308
rect 148410 128296 148416 128308
rect 147732 128268 148416 128296
rect 147732 128256 147738 128268
rect 148410 128256 148416 128268
rect 148468 128256 148474 128308
rect 232682 126896 232688 126948
rect 232740 126936 232746 126948
rect 239766 126936 239772 126948
rect 232740 126908 239772 126936
rect 232740 126896 232746 126908
rect 239766 126896 239772 126908
rect 239824 126896 239830 126948
rect 483658 126896 483664 126948
rect 483716 126936 483722 126948
rect 491662 126936 491668 126948
rect 483716 126908 491668 126936
rect 483716 126896 483722 126908
rect 491662 126896 491668 126908
rect 491720 126896 491726 126948
rect 512730 126896 512736 126948
rect 512788 126936 512794 126948
rect 519630 126936 519636 126948
rect 512788 126908 519636 126936
rect 512788 126896 512794 126908
rect 519630 126896 519636 126908
rect 519688 126896 519694 126948
rect 428642 126216 428648 126268
rect 428700 126256 428706 126268
rect 435726 126256 435732 126268
rect 428700 126228 435732 126256
rect 428700 126216 428706 126228
rect 435726 126216 435732 126228
rect 435784 126216 435790 126268
rect 287698 126080 287704 126132
rect 287756 126120 287762 126132
rect 295702 126120 295708 126132
rect 287756 126092 295708 126120
rect 287756 126080 287762 126092
rect 295702 126080 295708 126092
rect 295760 126080 295766 126132
rect 316770 126080 316776 126132
rect 316828 126120 316834 126132
rect 323670 126120 323676 126132
rect 316828 126092 323676 126120
rect 316828 126080 316834 126092
rect 323670 126080 323676 126092
rect 323728 126080 323734 126132
rect 13722 125536 13728 125588
rect 13780 125576 13786 125588
rect 66254 125576 66260 125588
rect 13780 125548 66260 125576
rect 13780 125536 13786 125548
rect 66254 125536 66260 125548
rect 66312 125536 66318 125588
rect 70302 125536 70308 125588
rect 70360 125576 70366 125588
rect 121454 125576 121460 125588
rect 70360 125548 121460 125576
rect 70360 125536 70366 125548
rect 121454 125536 121460 125548
rect 121512 125536 121518 125588
rect 126882 125536 126888 125588
rect 126940 125576 126946 125588
rect 178034 125576 178040 125588
rect 126940 125548 178040 125576
rect 126940 125536 126946 125548
rect 178034 125536 178040 125548
rect 178092 125536 178098 125588
rect 209682 125536 209688 125588
rect 209740 125576 209746 125588
rect 262214 125576 262220 125588
rect 209740 125548 262220 125576
rect 209740 125536 209746 125548
rect 262214 125536 262220 125548
rect 262272 125536 262278 125588
rect 266262 125536 266268 125588
rect 266320 125576 266326 125588
rect 317414 125576 317420 125588
rect 266320 125548 317420 125576
rect 266320 125536 266326 125548
rect 317414 125536 317420 125548
rect 317472 125536 317478 125588
rect 322842 125536 322848 125588
rect 322900 125576 322906 125588
rect 373994 125576 374000 125588
rect 322900 125548 374000 125576
rect 322900 125536 322906 125548
rect 373994 125536 374000 125548
rect 374052 125536 374058 125588
rect 405642 125536 405648 125588
rect 405700 125576 405706 125588
rect 458174 125576 458180 125588
rect 405700 125548 458180 125576
rect 405700 125536 405706 125548
rect 458174 125536 458180 125548
rect 458232 125536 458238 125588
rect 489822 125536 489828 125588
rect 489880 125576 489886 125588
rect 542354 125576 542360 125588
rect 489880 125548 542360 125576
rect 489880 125536 489886 125548
rect 542354 125536 542360 125548
rect 542412 125536 542418 125588
rect 42702 125468 42708 125520
rect 42760 125508 42766 125520
rect 93854 125508 93860 125520
rect 42760 125480 93860 125508
rect 42760 125468 42766 125480
rect 93854 125468 93860 125480
rect 93912 125468 93918 125520
rect 97902 125468 97908 125520
rect 97960 125508 97966 125520
rect 149054 125508 149060 125520
rect 97960 125480 149060 125508
rect 97960 125468 97966 125480
rect 149054 125468 149060 125480
rect 149112 125468 149118 125520
rect 154482 125468 154488 125520
rect 154540 125508 154546 125520
rect 205634 125508 205640 125520
rect 154540 125480 205640 125508
rect 154540 125468 154546 125480
rect 205634 125468 205640 125480
rect 205692 125468 205698 125520
rect 238662 125468 238668 125520
rect 238720 125508 238726 125520
rect 289814 125508 289820 125520
rect 238720 125480 289820 125508
rect 238720 125468 238726 125480
rect 289814 125468 289820 125480
rect 289872 125468 289878 125520
rect 293862 125468 293868 125520
rect 293920 125508 293926 125520
rect 345014 125508 345020 125520
rect 293920 125480 345020 125508
rect 293920 125468 293926 125480
rect 345014 125468 345020 125480
rect 345072 125468 345078 125520
rect 350442 125468 350448 125520
rect 350500 125508 350506 125520
rect 401594 125508 401600 125520
rect 350500 125480 401600 125508
rect 350500 125468 350506 125480
rect 401594 125468 401600 125480
rect 401652 125468 401658 125520
rect 434622 125468 434628 125520
rect 434680 125508 434686 125520
rect 485774 125508 485780 125520
rect 434680 125480 485780 125508
rect 434680 125468 434686 125480
rect 485774 125468 485780 125480
rect 485832 125468 485838 125520
rect 518802 125468 518808 125520
rect 518860 125508 518866 125520
rect 569954 125508 569960 125520
rect 518860 125480 569960 125508
rect 518860 125468 518866 125480
rect 569954 125468 569960 125480
rect 570012 125468 570018 125520
rect 182082 125400 182088 125452
rect 182140 125440 182146 125452
rect 233234 125440 233240 125452
rect 182140 125412 233240 125440
rect 182140 125400 182146 125412
rect 233234 125400 233240 125412
rect 233292 125400 233298 125452
rect 378042 125400 378048 125452
rect 378100 125440 378106 125452
rect 429194 125440 429200 125452
rect 378100 125412 429200 125440
rect 378100 125400 378106 125412
rect 429194 125400 429200 125412
rect 429252 125400 429258 125452
rect 462222 125400 462228 125452
rect 462280 125440 462286 125452
rect 513374 125440 513380 125452
rect 462280 125412 513380 125440
rect 462280 125400 462286 125412
rect 513374 125400 513380 125412
rect 513432 125400 513438 125452
rect 35618 124788 35624 124840
rect 35676 124828 35682 124840
rect 36906 124828 36912 124840
rect 35676 124800 36912 124828
rect 35676 124788 35682 124800
rect 36906 124788 36912 124800
rect 36964 124788 36970 124840
rect 343542 124788 343548 124840
rect 343600 124828 343606 124840
rect 345658 124828 345664 124840
rect 343600 124800 345664 124828
rect 343600 124788 343606 124800
rect 345658 124788 345664 124800
rect 345716 124788 345722 124840
rect 178678 122748 178684 122800
rect 178736 122788 178742 122800
rect 184014 122788 184020 122800
rect 178736 122760 184020 122788
rect 178736 122748 178742 122760
rect 184014 122748 184020 122760
rect 184072 122748 184078 122800
rect 231578 122748 231584 122800
rect 231636 122788 231642 122800
rect 232498 122788 232504 122800
rect 231636 122760 232504 122788
rect 231636 122748 231642 122760
rect 232498 122748 232504 122760
rect 232556 122748 232562 122800
rect 374638 122748 374644 122800
rect 374696 122788 374702 122800
rect 379698 122788 379704 122800
rect 374696 122760 379704 122788
rect 374696 122748 374702 122760
rect 379698 122748 379704 122760
rect 379756 122748 379762 122800
rect 539318 122748 539324 122800
rect 539376 122788 539382 122800
rect 542998 122788 543004 122800
rect 539376 122760 543004 122788
rect 539376 122748 539382 122760
rect 542998 122748 543004 122760
rect 543056 122748 543062 122800
rect 36814 122680 36820 122732
rect 36872 122720 36878 122732
rect 557534 122720 557540 122732
rect 36872 122692 557540 122720
rect 36872 122680 36878 122692
rect 557534 122680 557540 122692
rect 557592 122680 557598 122732
rect 15194 122612 15200 122664
rect 15252 122652 15258 122664
rect 43990 122652 43996 122664
rect 15252 122624 43996 122652
rect 15252 122612 15258 122624
rect 43990 122612 43996 122624
rect 44048 122612 44054 122664
rect 45526 122624 69796 122652
rect 25682 122544 25688 122596
rect 25740 122584 25746 122596
rect 36998 122584 37004 122596
rect 25740 122556 37004 122584
rect 25740 122544 25746 122556
rect 36998 122544 37004 122556
rect 37056 122544 37062 122596
rect 42886 122544 42892 122596
rect 42944 122584 42950 122596
rect 45526 122584 45554 122624
rect 42944 122556 45554 122584
rect 42944 122544 42950 122556
rect 53650 122544 53656 122596
rect 53708 122584 53714 122596
rect 69658 122584 69664 122596
rect 53708 122556 69664 122584
rect 53708 122544 53714 122556
rect 69658 122544 69664 122556
rect 69716 122544 69722 122596
rect 69768 122584 69796 122624
rect 71866 122612 71872 122664
rect 71924 122652 71930 122664
rect 100018 122652 100024 122664
rect 71924 122624 100024 122652
rect 71924 122612 71930 122624
rect 100018 122612 100024 122624
rect 100076 122612 100082 122664
rect 127986 122652 127992 122664
rect 103486 122624 127992 122652
rect 71958 122584 71964 122596
rect 69768 122556 71964 122584
rect 71958 122544 71964 122556
rect 72016 122544 72022 122596
rect 81986 122544 81992 122596
rect 82044 122584 82050 122596
rect 94498 122584 94504 122596
rect 82044 122556 94504 122584
rect 82044 122544 82050 122556
rect 94498 122544 94504 122556
rect 94556 122544 94562 122596
rect 99466 122544 99472 122596
rect 99524 122584 99530 122596
rect 103486 122584 103514 122624
rect 127986 122612 127992 122624
rect 128044 122612 128050 122664
rect 155954 122652 155960 122664
rect 132466 122624 155960 122652
rect 99524 122556 103514 122584
rect 99524 122544 99530 122556
rect 109678 122544 109684 122596
rect 109736 122584 109742 122596
rect 120718 122584 120724 122596
rect 109736 122556 120724 122584
rect 109736 122544 109742 122556
rect 120718 122544 120724 122556
rect 120776 122544 120782 122596
rect 127066 122544 127072 122596
rect 127124 122584 127130 122596
rect 132466 122584 132494 122624
rect 155954 122612 155960 122624
rect 156012 122612 156018 122664
rect 165982 122612 165988 122664
rect 166040 122652 166046 122664
rect 177298 122652 177304 122664
rect 166040 122624 177304 122652
rect 166040 122612 166046 122624
rect 177298 122612 177304 122624
rect 177356 122612 177362 122664
rect 183646 122612 183652 122664
rect 183704 122652 183710 122664
rect 211706 122652 211712 122664
rect 183704 122624 211712 122652
rect 183704 122612 183710 122624
rect 211706 122612 211712 122624
rect 211764 122612 211770 122664
rect 221918 122612 221924 122664
rect 221976 122652 221982 122664
rect 232590 122652 232596 122664
rect 221976 122624 232596 122652
rect 221976 122612 221982 122624
rect 232590 122612 232596 122624
rect 232648 122612 232654 122664
rect 238846 122612 238852 122664
rect 238904 122652 238910 122664
rect 268010 122652 268016 122664
rect 238904 122624 268016 122652
rect 238904 122612 238910 122624
rect 268010 122612 268016 122624
rect 268068 122612 268074 122664
rect 277670 122612 277676 122664
rect 277728 122652 277734 122664
rect 289078 122652 289084 122664
rect 277728 122624 289084 122652
rect 277728 122612 277734 122624
rect 289078 122612 289084 122624
rect 289136 122612 289142 122664
rect 306006 122612 306012 122664
rect 306064 122652 306070 122664
rect 316678 122652 316684 122664
rect 306064 122624 316684 122652
rect 306064 122612 306070 122624
rect 316678 122612 316684 122624
rect 316736 122612 316742 122664
rect 323026 122612 323032 122664
rect 323084 122652 323090 122664
rect 352006 122652 352012 122664
rect 323084 122624 352012 122652
rect 323084 122612 323090 122624
rect 352006 122612 352012 122624
rect 352064 122612 352070 122664
rect 361666 122612 361672 122664
rect 361724 122652 361730 122664
rect 373258 122652 373264 122664
rect 361724 122624 373264 122652
rect 361724 122612 361730 122624
rect 373258 122612 373264 122624
rect 373316 122612 373322 122664
rect 379606 122612 379612 122664
rect 379664 122652 379670 122664
rect 408034 122652 408040 122664
rect 379664 122624 408040 122652
rect 379664 122612 379670 122624
rect 408034 122612 408040 122624
rect 408092 122612 408098 122664
rect 417694 122612 417700 122664
rect 417752 122652 417758 122664
rect 428550 122652 428556 122664
rect 417752 122624 428556 122652
rect 417752 122612 417758 122624
rect 428550 122612 428556 122624
rect 428608 122612 428614 122664
rect 434806 122612 434812 122664
rect 434864 122652 434870 122664
rect 463786 122652 463792 122664
rect 434864 122624 463792 122652
rect 434864 122612 434870 122624
rect 463786 122612 463792 122624
rect 463844 122612 463850 122664
rect 473998 122612 474004 122664
rect 474056 122652 474062 122664
rect 485038 122652 485044 122664
rect 474056 122624 485044 122652
rect 474056 122612 474062 122624
rect 485038 122612 485044 122624
rect 485096 122612 485102 122664
rect 501690 122612 501696 122664
rect 501748 122652 501754 122664
rect 512638 122652 512644 122664
rect 501748 122624 512644 122652
rect 501748 122612 501754 122624
rect 512638 122612 512644 122624
rect 512696 122612 512702 122664
rect 518986 122612 518992 122664
rect 519044 122652 519050 122664
rect 547874 122652 547880 122664
rect 519044 122624 547880 122652
rect 519044 122612 519050 122624
rect 547874 122612 547880 122624
rect 547932 122612 547938 122664
rect 127124 122556 132494 122584
rect 127124 122544 127130 122556
rect 137646 122544 137652 122596
rect 137704 122584 137710 122596
rect 148318 122584 148324 122596
rect 137704 122556 148324 122584
rect 137704 122544 137710 122556
rect 148318 122544 148324 122556
rect 148376 122544 148382 122596
rect 193674 122544 193680 122596
rect 193732 122584 193738 122596
rect 204898 122584 204904 122596
rect 193732 122556 204904 122584
rect 193732 122544 193738 122556
rect 204898 122544 204904 122556
rect 204956 122544 204962 122596
rect 249702 122544 249708 122596
rect 249760 122584 249766 122596
rect 260190 122584 260196 122596
rect 249760 122556 260196 122584
rect 249760 122544 249766 122556
rect 260190 122544 260196 122556
rect 260248 122544 260254 122596
rect 333698 122544 333704 122596
rect 333756 122584 333762 122596
rect 344278 122584 344284 122596
rect 333756 122556 344284 122584
rect 333756 122544 333762 122556
rect 344278 122544 344284 122556
rect 344336 122544 344342 122596
rect 390002 122544 390008 122596
rect 390060 122584 390066 122596
rect 400858 122584 400864 122596
rect 390060 122556 400864 122584
rect 390060 122544 390066 122556
rect 400858 122544 400864 122556
rect 400916 122544 400922 122596
rect 445662 122544 445668 122596
rect 445720 122584 445726 122596
rect 456150 122584 456156 122596
rect 445720 122556 456156 122584
rect 445720 122544 445726 122556
rect 456150 122544 456156 122556
rect 456208 122544 456214 122596
rect 529658 122544 529664 122596
rect 529716 122584 529722 122596
rect 540238 122584 540244 122596
rect 529716 122556 540244 122584
rect 529716 122544 529722 122556
rect 540238 122544 540244 122556
rect 540296 122544 540302 122596
rect 39298 122476 39304 122528
rect 39356 122516 39362 122528
rect 567194 122516 567200 122528
rect 39356 122488 567200 122516
rect 39356 122476 39362 122488
rect 567194 122476 567200 122488
rect 567252 122476 567258 122528
rect 16022 119348 16028 119400
rect 16080 119388 16086 119400
rect 547874 119388 547880 119400
rect 16080 119360 547880 119388
rect 16080 119348 16086 119360
rect 547874 119348 547880 119360
rect 547932 119348 547938 119400
rect 25682 118940 25688 118992
rect 25740 118980 25746 118992
rect 261478 118980 261484 118992
rect 25740 118952 261484 118980
rect 25740 118940 25746 118952
rect 261478 118940 261484 118952
rect 261536 118940 261542 118992
rect 148318 118872 148324 118924
rect 148376 118912 148382 118924
rect 165706 118912 165712 118924
rect 148376 118884 165712 118912
rect 148376 118872 148382 118884
rect 165706 118872 165712 118884
rect 165764 118872 165770 118924
rect 175458 118872 175464 118924
rect 175516 118912 175522 118924
rect 193674 118912 193680 118924
rect 175516 118884 193680 118912
rect 175516 118872 175522 118884
rect 193674 118872 193680 118884
rect 193732 118872 193738 118924
rect 203518 118872 203524 118924
rect 203576 118912 203582 118924
rect 221366 118912 221372 118924
rect 203576 118884 221372 118912
rect 203576 118872 203582 118884
rect 221366 118872 221372 118884
rect 221424 118872 221430 118924
rect 408034 118872 408040 118924
rect 408092 118912 408098 118924
rect 428642 118912 428648 118924
rect 408092 118884 428648 118912
rect 408092 118872 408098 118884
rect 428642 118872 428648 118884
rect 428700 118872 428706 118924
rect 492030 118872 492036 118924
rect 492088 118912 492094 118924
rect 512730 118912 512736 118924
rect 492088 118884 512736 118912
rect 492088 118872 492094 118884
rect 512730 118872 512736 118884
rect 512788 118872 512794 118924
rect 36906 118804 36912 118856
rect 36964 118844 36970 118856
rect 53650 118844 53656 118856
rect 36964 118816 53656 118844
rect 36964 118804 36970 118816
rect 53650 118804 53656 118816
rect 53708 118804 53714 118856
rect 64322 118804 64328 118856
rect 64380 118844 64386 118856
rect 81434 118844 81440 118856
rect 64380 118816 81440 118844
rect 64380 118804 64386 118816
rect 81434 118804 81440 118816
rect 81492 118804 81498 118856
rect 91462 118804 91468 118856
rect 91520 118844 91526 118856
rect 109678 118844 109684 118856
rect 91520 118816 109684 118844
rect 91520 118804 91526 118816
rect 109678 118804 109684 118816
rect 109736 118804 109742 118856
rect 119430 118804 119436 118856
rect 119488 118844 119494 118856
rect 137646 118844 137652 118856
rect 119488 118816 137652 118844
rect 119488 118804 119494 118816
rect 137646 118804 137652 118816
rect 137704 118804 137710 118856
rect 156322 118804 156328 118856
rect 156380 118844 156386 118856
rect 178678 118844 178684 118856
rect 156380 118816 178684 118844
rect 156380 118804 156386 118816
rect 178678 118804 178684 118816
rect 178736 118804 178742 118856
rect 232590 118804 232596 118856
rect 232648 118844 232654 118856
rect 249702 118844 249708 118856
rect 232648 118816 249708 118844
rect 232648 118804 232654 118816
rect 249702 118804 249708 118816
rect 249760 118804 249766 118856
rect 260098 118804 260104 118856
rect 260156 118844 260162 118856
rect 277670 118844 277676 118856
rect 260156 118816 277676 118844
rect 260156 118804 260162 118816
rect 277670 118804 277676 118816
rect 277728 118804 277734 118856
rect 287514 118804 287520 118856
rect 287572 118844 287578 118856
rect 305362 118844 305368 118856
rect 287572 118816 305368 118844
rect 287572 118804 287578 118816
rect 305362 118804 305368 118816
rect 305420 118804 305426 118856
rect 315482 118804 315488 118856
rect 315540 118844 315546 118856
rect 333698 118844 333704 118856
rect 315540 118816 333704 118844
rect 315540 118804 315546 118816
rect 333698 118804 333704 118816
rect 333756 118804 333762 118856
rect 345658 118804 345664 118856
rect 345716 118844 345722 118856
rect 361666 118844 361672 118856
rect 345716 118816 361672 118844
rect 345716 118804 345722 118816
rect 361666 118804 361672 118816
rect 361724 118804 361730 118856
rect 371510 118804 371516 118856
rect 371568 118844 371574 118856
rect 389358 118844 389364 118856
rect 371568 118816 389364 118844
rect 371568 118804 371574 118816
rect 389358 118804 389364 118816
rect 389416 118804 389422 118856
rect 399478 118804 399484 118856
rect 399536 118844 399542 118856
rect 417694 118844 417700 118856
rect 399536 118816 417700 118844
rect 399536 118804 399542 118816
rect 417694 118804 417700 118816
rect 417752 118804 417758 118856
rect 456150 118804 456156 118856
rect 456208 118844 456214 118856
rect 473354 118844 473360 118856
rect 456208 118816 473360 118844
rect 456208 118804 456214 118816
rect 473354 118804 473360 118816
rect 473412 118804 473418 118856
rect 483474 118804 483480 118856
rect 483532 118844 483538 118856
rect 501690 118844 501696 118856
rect 483532 118816 501696 118844
rect 483532 118804 483538 118816
rect 501690 118804 501696 118816
rect 501748 118804 501754 118856
rect 36998 118736 37004 118788
rect 37056 118776 37062 118788
rect 63310 118776 63316 118788
rect 37056 118748 63316 118776
rect 37056 118736 37062 118748
rect 63310 118736 63316 118748
rect 63368 118736 63374 118788
rect 66898 118736 66904 118788
rect 66956 118776 66962 118788
rect 91094 118776 91100 118788
rect 66956 118748 91100 118776
rect 66956 118736 66962 118748
rect 91094 118736 91100 118748
rect 91152 118736 91158 118788
rect 94498 118736 94504 118788
rect 94556 118776 94562 118788
rect 119338 118776 119344 118788
rect 94556 118748 119344 118776
rect 94556 118736 94562 118748
rect 119338 118736 119344 118748
rect 119396 118736 119402 118788
rect 120718 118736 120724 118788
rect 120776 118776 120782 118788
rect 147306 118776 147312 118788
rect 120776 118748 147312 118776
rect 120776 118736 120782 118748
rect 147306 118736 147312 118748
rect 147364 118736 147370 118788
rect 148410 118736 148416 118788
rect 148468 118776 148474 118788
rect 175366 118776 175372 118788
rect 148468 118748 175372 118776
rect 148468 118736 148474 118748
rect 175366 118736 175372 118748
rect 175424 118736 175430 118788
rect 177298 118736 177304 118788
rect 177356 118776 177362 118788
rect 203334 118776 203340 118788
rect 177356 118748 203340 118776
rect 177356 118736 177362 118748
rect 203334 118736 203340 118748
rect 203392 118736 203398 118788
rect 204898 118736 204904 118788
rect 204956 118776 204962 118788
rect 231026 118776 231032 118788
rect 204956 118748 231032 118776
rect 204956 118736 204962 118748
rect 231026 118736 231032 118748
rect 231084 118736 231090 118788
rect 232498 118736 232504 118788
rect 232556 118776 232562 118788
rect 259362 118776 259368 118788
rect 232556 118748 259368 118776
rect 232556 118736 232562 118748
rect 259362 118736 259368 118748
rect 259420 118736 259426 118788
rect 268010 118736 268016 118788
rect 268068 118776 268074 118788
rect 287698 118776 287704 118788
rect 268068 118748 287704 118776
rect 268068 118736 268074 118748
rect 287698 118736 287704 118748
rect 287756 118736 287762 118788
rect 296346 118736 296352 118788
rect 296404 118776 296410 118788
rect 316770 118776 316776 118788
rect 296404 118748 316776 118776
rect 296404 118736 296410 118748
rect 316770 118736 316776 118748
rect 316828 118736 316834 118788
rect 352006 118736 352012 118788
rect 352064 118776 352070 118788
rect 374638 118776 374644 118788
rect 352064 118748 374644 118776
rect 352064 118736 352070 118748
rect 374638 118736 374644 118748
rect 374696 118736 374702 118788
rect 428458 118736 428464 118788
rect 428516 118776 428522 118788
rect 445662 118776 445668 118788
rect 428516 118748 445668 118776
rect 428516 118736 428522 118748
rect 445662 118736 445668 118748
rect 445720 118736 445726 118788
rect 464338 118736 464344 118788
rect 464396 118776 464402 118788
rect 483658 118776 483664 118788
rect 464396 118748 483664 118776
rect 464396 118736 464402 118748
rect 483658 118736 483664 118748
rect 483716 118736 483722 118788
rect 511442 118736 511448 118788
rect 511500 118776 511506 118788
rect 529658 118776 529664 118788
rect 511500 118748 529664 118776
rect 511500 118736 511506 118748
rect 529658 118736 529664 118748
rect 529716 118736 529722 118788
rect 542998 118736 543004 118788
rect 543056 118776 543062 118788
rect 557534 118776 557540 118788
rect 543056 118748 557540 118776
rect 543056 118736 543062 118748
rect 557534 118736 557540 118748
rect 557592 118736 557598 118788
rect 212350 118668 212356 118720
rect 212408 118708 212414 118720
rect 232682 118708 232688 118720
rect 212408 118680 232688 118708
rect 212408 118668 212414 118680
rect 232682 118668 232688 118680
rect 232740 118668 232746 118720
rect 260190 118668 260196 118720
rect 260248 118708 260254 118720
rect 287330 118708 287336 118720
rect 260248 118680 287336 118708
rect 260248 118668 260254 118680
rect 287330 118668 287336 118680
rect 287388 118668 287394 118720
rect 289078 118668 289084 118720
rect 289136 118708 289142 118720
rect 315022 118708 315028 118720
rect 289136 118680 315028 118708
rect 289136 118668 289142 118680
rect 315022 118668 315028 118680
rect 315080 118668 315086 118720
rect 316678 118668 316684 118720
rect 316736 118708 316742 118720
rect 343358 118708 343364 118720
rect 316736 118680 343364 118708
rect 316736 118668 316742 118680
rect 343358 118668 343364 118680
rect 343416 118668 343422 118720
rect 344278 118668 344284 118720
rect 344336 118708 344342 118720
rect 371326 118708 371332 118720
rect 344336 118680 371332 118708
rect 344336 118668 344342 118680
rect 371326 118668 371332 118680
rect 371384 118668 371390 118720
rect 373258 118668 373264 118720
rect 373316 118708 373322 118720
rect 399018 118708 399024 118720
rect 373316 118680 399024 118708
rect 373316 118668 373322 118680
rect 399018 118668 399024 118680
rect 399076 118668 399082 118720
rect 400858 118668 400864 118720
rect 400916 118708 400922 118720
rect 427354 118708 427360 118720
rect 400916 118680 427360 118708
rect 400916 118668 400922 118680
rect 427354 118668 427360 118680
rect 427412 118668 427418 118720
rect 428550 118668 428556 118720
rect 428608 118708 428614 118720
rect 455322 118708 455328 118720
rect 428608 118680 455328 118708
rect 428608 118668 428614 118680
rect 455322 118668 455328 118680
rect 455380 118668 455386 118720
rect 456058 118668 456064 118720
rect 456116 118708 456122 118720
rect 483014 118708 483020 118720
rect 456116 118680 483020 118708
rect 456116 118668 456122 118680
rect 483014 118668 483020 118680
rect 483072 118668 483078 118720
rect 485038 118668 485044 118720
rect 485096 118708 485102 118720
rect 511350 118708 511356 118720
rect 485096 118680 511356 118708
rect 485096 118668 485102 118680
rect 511350 118668 511356 118680
rect 511408 118668 511414 118720
rect 512638 118668 512644 118720
rect 512696 118708 512702 118720
rect 539318 118708 539324 118720
rect 512696 118680 539324 118708
rect 512696 118668 512702 118680
rect 539318 118668 539324 118680
rect 539376 118668 539382 118720
rect 540238 118668 540244 118720
rect 540296 118708 540302 118720
rect 567194 118708 567200 118720
rect 540296 118680 567200 118708
rect 540296 118668 540302 118680
rect 567194 118668 567200 118680
rect 567252 118668 567258 118720
rect 37918 116560 37924 116612
rect 37976 116600 37982 116612
rect 545758 116600 545764 116612
rect 37976 116572 545764 116600
rect 37976 116560 37982 116572
rect 545758 116560 545764 116572
rect 545816 116560 545822 116612
rect 35618 116084 35624 116136
rect 35676 116124 35682 116136
rect 36814 116124 36820 116136
rect 35676 116096 36820 116124
rect 35676 116084 35682 116096
rect 36814 116084 36820 116096
rect 36872 116084 36878 116136
rect 63586 100240 63592 100292
rect 63644 100280 63650 100292
rect 64322 100280 64328 100292
rect 63644 100252 64328 100280
rect 63644 100240 63650 100252
rect 64322 100240 64328 100252
rect 64380 100240 64386 100292
rect 455690 100240 455696 100292
rect 455748 100280 455754 100292
rect 456150 100280 456156 100292
rect 455748 100252 456156 100280
rect 455748 100240 455754 100252
rect 456150 100240 456156 100252
rect 456208 100240 456214 100292
rect 316770 98880 316776 98932
rect 316828 98920 316834 98932
rect 323670 98920 323676 98932
rect 316828 98892 323676 98920
rect 316828 98880 316834 98892
rect 323670 98880 323676 98892
rect 323728 98880 323734 98932
rect 287698 98744 287704 98796
rect 287756 98784 287762 98796
rect 295702 98784 295708 98796
rect 287756 98756 295708 98784
rect 287756 98744 287762 98756
rect 295702 98744 295708 98756
rect 295760 98744 295766 98796
rect 428642 98608 428648 98660
rect 428700 98648 428706 98660
rect 435726 98648 435732 98660
rect 428700 98620 435732 98648
rect 428700 98608 428706 98620
rect 435726 98608 435732 98620
rect 435784 98608 435790 98660
rect 483658 98608 483664 98660
rect 483716 98648 483722 98660
rect 491662 98648 491668 98660
rect 483716 98620 491668 98648
rect 483716 98608 483722 98620
rect 491662 98608 491668 98620
rect 491720 98608 491726 98660
rect 512730 98540 512736 98592
rect 512788 98580 512794 98592
rect 519630 98580 519636 98592
rect 512788 98552 519636 98580
rect 512788 98540 512794 98552
rect 519630 98540 519636 98552
rect 519688 98540 519694 98592
rect 232682 98200 232688 98252
rect 232740 98240 232746 98252
rect 239766 98240 239772 98252
rect 232740 98212 239772 98240
rect 232740 98200 232746 98212
rect 239766 98200 239772 98212
rect 239824 98200 239830 98252
rect 13722 97928 13728 97980
rect 13780 97968 13786 97980
rect 66254 97968 66260 97980
rect 13780 97940 66260 97968
rect 13780 97928 13786 97940
rect 66254 97928 66260 97940
rect 66312 97928 66318 97980
rect 97902 97928 97908 97980
rect 97960 97968 97966 97980
rect 149054 97968 149060 97980
rect 97960 97940 149060 97968
rect 97960 97928 97966 97940
rect 149054 97928 149060 97940
rect 149112 97928 149118 97980
rect 154482 97928 154488 97980
rect 154540 97968 154546 97980
rect 205634 97968 205640 97980
rect 154540 97940 205640 97968
rect 154540 97928 154546 97940
rect 205634 97928 205640 97940
rect 205692 97928 205698 97980
rect 209682 97928 209688 97980
rect 209740 97968 209746 97980
rect 262214 97968 262220 97980
rect 209740 97940 262220 97968
rect 209740 97928 209746 97940
rect 262214 97928 262220 97940
rect 262272 97928 262278 97980
rect 266262 97928 266268 97980
rect 266320 97968 266326 97980
rect 317414 97968 317420 97980
rect 266320 97940 317420 97968
rect 266320 97928 266326 97940
rect 317414 97928 317420 97940
rect 317472 97928 317478 97980
rect 322842 97928 322848 97980
rect 322900 97968 322906 97980
rect 373994 97968 374000 97980
rect 322900 97940 374000 97968
rect 322900 97928 322906 97940
rect 373994 97928 374000 97940
rect 374052 97928 374058 97980
rect 405642 97928 405648 97980
rect 405700 97968 405706 97980
rect 458174 97968 458180 97980
rect 405700 97940 458180 97968
rect 405700 97928 405706 97940
rect 458174 97928 458180 97940
rect 458232 97928 458238 97980
rect 489822 97928 489828 97980
rect 489880 97968 489886 97980
rect 542354 97968 542360 97980
rect 489880 97940 542360 97968
rect 489880 97928 489886 97940
rect 542354 97928 542360 97940
rect 542412 97928 542418 97980
rect 42702 97860 42708 97912
rect 42760 97900 42766 97912
rect 93854 97900 93860 97912
rect 42760 97872 93860 97900
rect 42760 97860 42766 97872
rect 93854 97860 93860 97872
rect 93912 97860 93918 97912
rect 126882 97860 126888 97912
rect 126940 97900 126946 97912
rect 178034 97900 178040 97912
rect 126940 97872 178040 97900
rect 126940 97860 126946 97872
rect 178034 97860 178040 97872
rect 178092 97860 178098 97912
rect 182082 97860 182088 97912
rect 182140 97900 182146 97912
rect 233234 97900 233240 97912
rect 182140 97872 233240 97900
rect 182140 97860 182146 97872
rect 233234 97860 233240 97872
rect 233292 97860 233298 97912
rect 238662 97860 238668 97912
rect 238720 97900 238726 97912
rect 289814 97900 289820 97912
rect 238720 97872 289820 97900
rect 238720 97860 238726 97872
rect 289814 97860 289820 97872
rect 289872 97860 289878 97912
rect 293862 97860 293868 97912
rect 293920 97900 293926 97912
rect 345014 97900 345020 97912
rect 293920 97872 345020 97900
rect 293920 97860 293926 97872
rect 345014 97860 345020 97872
rect 345072 97860 345078 97912
rect 378042 97860 378048 97912
rect 378100 97900 378106 97912
rect 429194 97900 429200 97912
rect 378100 97872 429200 97900
rect 378100 97860 378106 97872
rect 429194 97860 429200 97872
rect 429252 97860 429258 97912
rect 462222 97860 462228 97912
rect 462280 97900 462286 97912
rect 513374 97900 513380 97912
rect 462280 97872 513380 97900
rect 462280 97860 462286 97872
rect 513374 97860 513380 97872
rect 513432 97860 513438 97912
rect 518802 97860 518808 97912
rect 518860 97900 518866 97912
rect 569954 97900 569960 97912
rect 518860 97872 569960 97900
rect 518860 97860 518866 97872
rect 569954 97860 569960 97872
rect 570012 97860 570018 97912
rect 70302 97792 70308 97844
rect 70360 97832 70366 97844
rect 121454 97832 121460 97844
rect 70360 97804 121460 97832
rect 70360 97792 70366 97804
rect 121454 97792 121460 97804
rect 121512 97792 121518 97844
rect 231670 97792 231676 97844
rect 231728 97832 231734 97844
rect 232590 97832 232596 97844
rect 231728 97804 232596 97832
rect 231728 97792 231734 97804
rect 232590 97792 232596 97804
rect 232648 97792 232654 97844
rect 350442 97792 350448 97844
rect 350500 97832 350506 97844
rect 401594 97832 401600 97844
rect 350500 97804 401600 97832
rect 350500 97792 350506 97804
rect 401594 97792 401600 97804
rect 401652 97792 401658 97844
rect 434622 97792 434628 97844
rect 434680 97832 434686 97844
rect 485774 97832 485780 97844
rect 434680 97804 485780 97832
rect 434680 97792 434686 97804
rect 485774 97792 485780 97804
rect 485832 97792 485838 97844
rect 539502 97792 539508 97844
rect 539560 97832 539566 97844
rect 542998 97832 543004 97844
rect 539560 97804 543004 97832
rect 539560 97792 539566 97804
rect 542998 97792 543004 97804
rect 543056 97792 543062 97844
rect 35618 97656 35624 97708
rect 35676 97696 35682 97708
rect 36906 97696 36912 97708
rect 35676 97668 36912 97696
rect 35676 97656 35682 97668
rect 36906 97656 36912 97668
rect 36964 97656 36970 97708
rect 343634 97656 343640 97708
rect 343692 97696 343698 97708
rect 345658 97696 345664 97708
rect 343692 97668 345664 97696
rect 343692 97656 343698 97668
rect 345658 97656 345664 97668
rect 345716 97656 345722 97708
rect 178678 95140 178684 95192
rect 178736 95180 178742 95192
rect 184014 95180 184020 95192
rect 178736 95152 184020 95180
rect 178736 95140 178742 95152
rect 184014 95140 184020 95152
rect 184072 95140 184078 95192
rect 374638 95140 374644 95192
rect 374696 95180 374702 95192
rect 379698 95180 379704 95192
rect 374696 95152 379704 95180
rect 374696 95140 374702 95152
rect 379698 95140 379704 95152
rect 379756 95140 379762 95192
rect 15194 95072 15200 95124
rect 15252 95112 15258 95124
rect 43990 95112 43996 95124
rect 15252 95084 43996 95112
rect 15252 95072 15258 95084
rect 43990 95072 43996 95084
rect 44048 95072 44054 95124
rect 71038 95072 71044 95124
rect 71096 95112 71102 95124
rect 567194 95112 567200 95124
rect 71096 95084 567200 95112
rect 71096 95072 71102 95084
rect 567194 95072 567200 95084
rect 567252 95072 567258 95124
rect 25682 95004 25688 95056
rect 25740 95044 25746 95056
rect 36998 95044 37004 95056
rect 25740 95016 37004 95044
rect 25740 95004 25746 95016
rect 36998 95004 37004 95016
rect 37056 95004 37062 95056
rect 53650 95004 53656 95056
rect 53708 95044 53714 95056
rect 66898 95044 66904 95056
rect 53708 95016 66904 95044
rect 53708 95004 53714 95016
rect 66898 95004 66904 95016
rect 66956 95004 66962 95056
rect 71866 95004 71872 95056
rect 71924 95044 71930 95056
rect 100018 95044 100024 95056
rect 71924 95016 100024 95044
rect 71924 95004 71930 95016
rect 100018 95004 100024 95016
rect 100076 95004 100082 95056
rect 127986 95044 127992 95056
rect 103486 95016 127992 95044
rect 42886 94936 42892 94988
rect 42944 94976 42950 94988
rect 72050 94976 72056 94988
rect 42944 94948 72056 94976
rect 42944 94936 42950 94948
rect 72050 94936 72056 94948
rect 72108 94936 72114 94988
rect 81986 94936 81992 94988
rect 82044 94976 82050 94988
rect 94498 94976 94504 94988
rect 82044 94948 94504 94976
rect 82044 94936 82050 94948
rect 94498 94936 94504 94948
rect 94556 94936 94562 94988
rect 99466 94936 99472 94988
rect 99524 94976 99530 94988
rect 103486 94976 103514 95016
rect 127986 95004 127992 95016
rect 128044 95004 128050 95056
rect 156046 95044 156052 95056
rect 132466 95016 156052 95044
rect 99524 94948 103514 94976
rect 99524 94936 99530 94948
rect 109678 94936 109684 94988
rect 109736 94976 109742 94988
rect 120718 94976 120724 94988
rect 109736 94948 120724 94976
rect 109736 94936 109742 94948
rect 120718 94936 120724 94948
rect 120776 94936 120782 94988
rect 127066 94936 127072 94988
rect 127124 94976 127130 94988
rect 132466 94976 132494 95016
rect 156046 95004 156052 95016
rect 156104 95004 156110 95056
rect 165982 95004 165988 95056
rect 166040 95044 166046 95056
rect 177298 95044 177304 95056
rect 166040 95016 177304 95044
rect 166040 95004 166046 95016
rect 177298 95004 177304 95016
rect 177356 95004 177362 95056
rect 183646 95004 183652 95056
rect 183704 95044 183710 95056
rect 211706 95044 211712 95056
rect 183704 95016 211712 95044
rect 183704 95004 183710 95016
rect 211706 95004 211712 95016
rect 211764 95004 211770 95056
rect 222010 95004 222016 95056
rect 222068 95044 222074 95056
rect 232498 95044 232504 95056
rect 222068 95016 232504 95044
rect 222068 95004 222074 95016
rect 232498 95004 232504 95016
rect 232556 95004 232562 95056
rect 238846 95004 238852 95056
rect 238904 95044 238910 95056
rect 268010 95044 268016 95056
rect 238904 95016 268016 95044
rect 238904 95004 238910 95016
rect 268010 95004 268016 95016
rect 268068 95004 268074 95056
rect 277670 95004 277676 95056
rect 277728 95044 277734 95056
rect 289078 95044 289084 95056
rect 277728 95016 289084 95044
rect 277728 95004 277734 95016
rect 289078 95004 289084 95016
rect 289136 95004 289142 95056
rect 306006 95004 306012 95056
rect 306064 95044 306070 95056
rect 316678 95044 316684 95056
rect 306064 95016 316684 95044
rect 306064 95004 306070 95016
rect 316678 95004 316684 95016
rect 316736 95004 316742 95056
rect 323026 95004 323032 95056
rect 323084 95044 323090 95056
rect 352006 95044 352012 95056
rect 323084 95016 352012 95044
rect 323084 95004 323090 95016
rect 352006 95004 352012 95016
rect 352064 95004 352070 95056
rect 361666 95004 361672 95056
rect 361724 95044 361730 95056
rect 373258 95044 373264 95056
rect 361724 95016 373264 95044
rect 361724 95004 361730 95016
rect 373258 95004 373264 95016
rect 373316 95004 373322 95056
rect 379606 95004 379612 95056
rect 379664 95044 379670 95056
rect 408034 95044 408040 95056
rect 379664 95016 408040 95044
rect 379664 95004 379670 95016
rect 408034 95004 408040 95016
rect 408092 95004 408098 95056
rect 417694 95004 417700 95056
rect 417752 95044 417758 95056
rect 428550 95044 428556 95056
rect 417752 95016 428556 95044
rect 417752 95004 417758 95016
rect 428550 95004 428556 95016
rect 428608 95004 428614 95056
rect 434806 95004 434812 95056
rect 434864 95044 434870 95056
rect 463694 95044 463700 95056
rect 434864 95016 463700 95044
rect 434864 95004 434870 95016
rect 463694 95004 463700 95016
rect 463752 95004 463758 95056
rect 473998 95004 474004 95056
rect 474056 95044 474062 95056
rect 485038 95044 485044 95056
rect 474056 95016 485044 95044
rect 474056 95004 474062 95016
rect 485038 95004 485044 95016
rect 485096 95004 485102 95056
rect 501690 95004 501696 95056
rect 501748 95044 501754 95056
rect 512638 95044 512644 95056
rect 501748 95016 512644 95044
rect 501748 95004 501754 95016
rect 512638 95004 512644 95016
rect 512696 95004 512702 95056
rect 518986 95004 518992 95056
rect 519044 95044 519050 95056
rect 547874 95044 547880 95056
rect 519044 95016 547880 95044
rect 519044 95004 519050 95016
rect 547874 95004 547880 95016
rect 547932 95004 547938 95056
rect 127124 94948 132494 94976
rect 127124 94936 127130 94948
rect 137646 94936 137652 94988
rect 137704 94976 137710 94988
rect 148410 94976 148416 94988
rect 137704 94948 148416 94976
rect 137704 94936 137710 94948
rect 148410 94936 148416 94948
rect 148468 94936 148474 94988
rect 193674 94936 193680 94988
rect 193732 94976 193738 94988
rect 204898 94976 204904 94988
rect 193732 94948 204904 94976
rect 193732 94936 193738 94948
rect 204898 94936 204904 94948
rect 204956 94936 204962 94988
rect 249702 94936 249708 94988
rect 249760 94976 249766 94988
rect 260190 94976 260196 94988
rect 249760 94948 260196 94976
rect 249760 94936 249766 94948
rect 260190 94936 260196 94948
rect 260248 94936 260254 94988
rect 333698 94936 333704 94988
rect 333756 94976 333762 94988
rect 344278 94976 344284 94988
rect 333756 94948 344284 94976
rect 333756 94936 333762 94948
rect 344278 94936 344284 94948
rect 344336 94936 344342 94988
rect 390002 94936 390008 94988
rect 390060 94976 390066 94988
rect 400858 94976 400864 94988
rect 390060 94948 400864 94976
rect 390060 94936 390066 94948
rect 400858 94936 400864 94948
rect 400916 94936 400922 94988
rect 445662 94936 445668 94988
rect 445720 94976 445726 94988
rect 456058 94976 456064 94988
rect 445720 94948 456064 94976
rect 445720 94936 445726 94948
rect 456058 94936 456064 94948
rect 456116 94936 456122 94988
rect 529658 94936 529664 94988
rect 529716 94976 529722 94988
rect 540238 94976 540244 94988
rect 529716 94948 540244 94976
rect 529716 94936 529722 94948
rect 540238 94936 540244 94948
rect 540296 94936 540302 94988
rect 36722 94868 36728 94920
rect 36780 94908 36786 94920
rect 557534 94908 557540 94920
rect 36780 94880 557540 94908
rect 36780 94868 36786 94880
rect 557534 94868 557540 94880
rect 557592 94868 557598 94920
rect 15286 91740 15292 91792
rect 15344 91780 15350 91792
rect 547874 91780 547880 91792
rect 15344 91752 547880 91780
rect 15344 91740 15350 91752
rect 547874 91740 547880 91752
rect 547932 91740 547938 91792
rect 25682 91264 25688 91316
rect 25740 91304 25746 91316
rect 71038 91304 71044 91316
rect 25740 91276 71044 91304
rect 25740 91264 25746 91276
rect 71038 91264 71044 91276
rect 71096 91264 71102 91316
rect 212350 91264 212356 91316
rect 212408 91304 212414 91316
rect 232682 91304 232688 91316
rect 212408 91276 232688 91304
rect 212408 91264 212414 91276
rect 232682 91264 232688 91276
rect 232740 91264 232746 91316
rect 296346 91264 296352 91316
rect 296404 91304 296410 91316
rect 316770 91304 316776 91316
rect 296404 91276 316776 91304
rect 296404 91264 296410 91276
rect 316770 91264 316776 91276
rect 316828 91264 316834 91316
rect 408034 91264 408040 91316
rect 408092 91304 408098 91316
rect 428642 91304 428648 91316
rect 408092 91276 428648 91304
rect 408092 91264 408098 91276
rect 428642 91264 428648 91276
rect 428700 91264 428706 91316
rect 36906 91196 36912 91248
rect 36964 91236 36970 91248
rect 53650 91236 53656 91248
rect 36964 91208 53656 91236
rect 36964 91196 36970 91208
rect 53650 91196 53656 91208
rect 53708 91196 53714 91248
rect 148318 91196 148324 91248
rect 148376 91236 148382 91248
rect 165706 91236 165712 91248
rect 148376 91208 165712 91236
rect 148376 91196 148382 91208
rect 165706 91196 165712 91208
rect 165764 91196 165770 91248
rect 175458 91196 175464 91248
rect 175516 91236 175522 91248
rect 193674 91236 193680 91248
rect 175516 91208 193680 91236
rect 175516 91196 175522 91208
rect 193674 91196 193680 91208
rect 193732 91196 193738 91248
rect 203518 91196 203524 91248
rect 203576 91236 203582 91248
rect 221366 91236 221372 91248
rect 203576 91208 221372 91236
rect 203576 91196 203582 91208
rect 221366 91196 221372 91208
rect 221424 91196 221430 91248
rect 260190 91196 260196 91248
rect 260248 91236 260254 91248
rect 277670 91236 277676 91248
rect 260248 91208 277676 91236
rect 260248 91196 260254 91208
rect 277670 91196 277676 91208
rect 277728 91196 277734 91248
rect 287514 91196 287520 91248
rect 287572 91236 287578 91248
rect 305362 91236 305368 91248
rect 287572 91208 305368 91236
rect 287572 91196 287578 91208
rect 305362 91196 305368 91208
rect 305420 91196 305426 91248
rect 345658 91196 345664 91248
rect 345716 91236 345722 91248
rect 361666 91236 361672 91248
rect 345716 91208 361672 91236
rect 345716 91196 345722 91208
rect 361666 91196 361672 91208
rect 361724 91196 361730 91248
rect 371510 91196 371516 91248
rect 371568 91236 371574 91248
rect 389358 91236 389364 91248
rect 371568 91208 389364 91236
rect 371568 91196 371574 91208
rect 389358 91196 389364 91208
rect 389416 91196 389422 91248
rect 399478 91196 399484 91248
rect 399536 91236 399542 91248
rect 417694 91236 417700 91248
rect 399536 91208 417700 91236
rect 399536 91196 399542 91208
rect 417694 91196 417700 91208
rect 417752 91196 417758 91248
rect 456150 91196 456156 91248
rect 456208 91236 456214 91248
rect 473354 91236 473360 91248
rect 456208 91208 473360 91236
rect 456208 91196 456214 91208
rect 473354 91196 473360 91208
rect 473412 91196 473418 91248
rect 483474 91196 483480 91248
rect 483532 91236 483538 91248
rect 501690 91236 501696 91248
rect 483532 91208 501696 91236
rect 483532 91196 483538 91208
rect 501690 91196 501696 91208
rect 501748 91196 501754 91248
rect 511442 91196 511448 91248
rect 511500 91236 511506 91248
rect 529658 91236 529664 91248
rect 511500 91208 529664 91236
rect 511500 91196 511506 91208
rect 529658 91196 529664 91208
rect 529716 91196 529722 91248
rect 36998 91128 37004 91180
rect 37056 91168 37062 91180
rect 63310 91168 63316 91180
rect 37056 91140 63316 91168
rect 37056 91128 37062 91140
rect 63310 91128 63316 91140
rect 63368 91128 63374 91180
rect 64322 91128 64328 91180
rect 64380 91168 64386 91180
rect 81434 91168 81440 91180
rect 64380 91140 81440 91168
rect 64380 91128 64386 91140
rect 81434 91128 81440 91140
rect 81492 91128 81498 91180
rect 91462 91128 91468 91180
rect 91520 91168 91526 91180
rect 109678 91168 109684 91180
rect 91520 91140 109684 91168
rect 91520 91128 91526 91140
rect 109678 91128 109684 91140
rect 109736 91128 109742 91180
rect 119430 91128 119436 91180
rect 119488 91168 119494 91180
rect 137646 91168 137652 91180
rect 119488 91140 137652 91168
rect 119488 91128 119494 91140
rect 137646 91128 137652 91140
rect 137704 91128 137710 91180
rect 156322 91128 156328 91180
rect 156380 91168 156386 91180
rect 178678 91168 178684 91180
rect 156380 91140 178684 91168
rect 156380 91128 156386 91140
rect 178678 91128 178684 91140
rect 178736 91128 178742 91180
rect 232590 91128 232596 91180
rect 232648 91168 232654 91180
rect 249702 91168 249708 91180
rect 232648 91140 249708 91168
rect 232648 91128 232654 91140
rect 249702 91128 249708 91140
rect 249760 91128 249766 91180
rect 268010 91128 268016 91180
rect 268068 91168 268074 91180
rect 287698 91168 287704 91180
rect 268068 91140 287704 91168
rect 268068 91128 268074 91140
rect 287698 91128 287704 91140
rect 287756 91128 287762 91180
rect 315482 91128 315488 91180
rect 315540 91168 315546 91180
rect 333698 91168 333704 91180
rect 315540 91140 333704 91168
rect 315540 91128 315546 91140
rect 333698 91128 333704 91140
rect 333756 91128 333762 91180
rect 352006 91128 352012 91180
rect 352064 91168 352070 91180
rect 374638 91168 374644 91180
rect 352064 91140 374644 91168
rect 352064 91128 352070 91140
rect 374638 91128 374644 91140
rect 374696 91128 374702 91180
rect 428458 91128 428464 91180
rect 428516 91168 428522 91180
rect 445662 91168 445668 91180
rect 428516 91140 445668 91168
rect 428516 91128 428522 91140
rect 445662 91128 445668 91140
rect 445720 91128 445726 91180
rect 464338 91128 464344 91180
rect 464396 91168 464402 91180
rect 483658 91168 483664 91180
rect 464396 91140 483664 91168
rect 464396 91128 464402 91140
rect 483658 91128 483664 91140
rect 483716 91128 483722 91180
rect 492030 91128 492036 91180
rect 492088 91168 492094 91180
rect 512730 91168 512736 91180
rect 492088 91140 512736 91168
rect 492088 91128 492094 91140
rect 512730 91128 512736 91140
rect 512788 91128 512794 91180
rect 542998 91128 543004 91180
rect 543056 91168 543062 91180
rect 557534 91168 557540 91180
rect 543056 91140 557540 91168
rect 543056 91128 543062 91140
rect 557534 91128 557540 91140
rect 557592 91128 557598 91180
rect 69658 91060 69664 91112
rect 69716 91100 69722 91112
rect 91094 91100 91100 91112
rect 69716 91072 91100 91100
rect 69716 91060 69722 91072
rect 91094 91060 91100 91072
rect 91152 91060 91158 91112
rect 94498 91060 94504 91112
rect 94556 91100 94562 91112
rect 119338 91100 119344 91112
rect 94556 91072 119344 91100
rect 94556 91060 94562 91072
rect 119338 91060 119344 91072
rect 119396 91060 119402 91112
rect 120718 91060 120724 91112
rect 120776 91100 120782 91112
rect 147306 91100 147312 91112
rect 120776 91072 147312 91100
rect 120776 91060 120782 91072
rect 147306 91060 147312 91072
rect 147364 91060 147370 91112
rect 148410 91060 148416 91112
rect 148468 91100 148474 91112
rect 175366 91100 175372 91112
rect 148468 91072 175372 91100
rect 148468 91060 148474 91072
rect 175366 91060 175372 91072
rect 175424 91060 175430 91112
rect 177298 91060 177304 91112
rect 177356 91100 177362 91112
rect 203334 91100 203340 91112
rect 177356 91072 203340 91100
rect 177356 91060 177362 91072
rect 203334 91060 203340 91072
rect 203392 91060 203398 91112
rect 204898 91060 204904 91112
rect 204956 91100 204962 91112
rect 231026 91100 231032 91112
rect 204956 91072 231032 91100
rect 204956 91060 204962 91072
rect 231026 91060 231032 91072
rect 231084 91060 231090 91112
rect 232498 91060 232504 91112
rect 232556 91100 232562 91112
rect 259362 91100 259368 91112
rect 232556 91072 259368 91100
rect 232556 91060 232562 91072
rect 259362 91060 259368 91072
rect 259420 91060 259426 91112
rect 260098 91060 260104 91112
rect 260156 91100 260162 91112
rect 287330 91100 287336 91112
rect 260156 91072 287336 91100
rect 260156 91060 260162 91072
rect 287330 91060 287336 91072
rect 287388 91060 287394 91112
rect 289078 91060 289084 91112
rect 289136 91100 289142 91112
rect 315022 91100 315028 91112
rect 289136 91072 315028 91100
rect 289136 91060 289142 91072
rect 315022 91060 315028 91072
rect 315080 91060 315086 91112
rect 316678 91060 316684 91112
rect 316736 91100 316742 91112
rect 343358 91100 343364 91112
rect 316736 91072 343364 91100
rect 316736 91060 316742 91072
rect 343358 91060 343364 91072
rect 343416 91060 343422 91112
rect 344278 91060 344284 91112
rect 344336 91100 344342 91112
rect 371326 91100 371332 91112
rect 344336 91072 371332 91100
rect 344336 91060 344342 91072
rect 371326 91060 371332 91072
rect 371384 91060 371390 91112
rect 373258 91060 373264 91112
rect 373316 91100 373322 91112
rect 399018 91100 399024 91112
rect 373316 91072 399024 91100
rect 373316 91060 373322 91072
rect 399018 91060 399024 91072
rect 399076 91060 399082 91112
rect 400858 91060 400864 91112
rect 400916 91100 400922 91112
rect 427354 91100 427360 91112
rect 400916 91072 427360 91100
rect 400916 91060 400922 91072
rect 427354 91060 427360 91072
rect 427412 91060 427418 91112
rect 428550 91060 428556 91112
rect 428608 91100 428614 91112
rect 455322 91100 455328 91112
rect 428608 91072 455328 91100
rect 428608 91060 428614 91072
rect 455322 91060 455328 91072
rect 455380 91060 455386 91112
rect 456058 91060 456064 91112
rect 456116 91100 456122 91112
rect 483014 91100 483020 91112
rect 456116 91072 483020 91100
rect 456116 91060 456122 91072
rect 483014 91060 483020 91072
rect 483072 91060 483078 91112
rect 485038 91060 485044 91112
rect 485096 91100 485102 91112
rect 511350 91100 511356 91112
rect 485096 91072 511356 91100
rect 485096 91060 485102 91072
rect 511350 91060 511356 91072
rect 511408 91060 511414 91112
rect 512638 91060 512644 91112
rect 512696 91100 512702 91112
rect 539318 91100 539324 91112
rect 512696 91072 539324 91100
rect 512696 91060 512702 91072
rect 539318 91060 539324 91072
rect 539376 91060 539382 91112
rect 540238 91060 540244 91112
rect 540296 91100 540302 91112
rect 567194 91100 567200 91112
rect 540296 91072 567200 91100
rect 540296 91060 540302 91072
rect 567194 91060 567200 91072
rect 567252 91060 567258 91112
rect 37918 90312 37924 90364
rect 37976 90352 37982 90364
rect 545758 90352 545764 90364
rect 37976 90324 545764 90352
rect 37976 90312 37982 90324
rect 545758 90312 545764 90324
rect 545816 90312 545822 90364
rect 35618 88408 35624 88460
rect 35676 88448 35682 88460
rect 36722 88448 36728 88460
rect 35676 88420 36728 88448
rect 35676 88408 35682 88420
rect 36722 88408 36728 88420
rect 36780 88408 36786 88460
rect 42702 88408 42708 88460
rect 42760 88448 42766 88460
rect 93854 88448 93860 88460
rect 42760 88420 93860 88448
rect 42760 88408 42766 88420
rect 93854 88408 93860 88420
rect 93912 88408 93918 88460
rect 154482 88408 154488 88460
rect 154540 88448 154546 88460
rect 205634 88448 205640 88460
rect 154540 88420 205640 88448
rect 154540 88408 154546 88420
rect 205634 88408 205640 88420
rect 205692 88408 205698 88460
rect 238662 88408 238668 88460
rect 238720 88448 238726 88460
rect 289814 88448 289820 88460
rect 238720 88420 289820 88448
rect 238720 88408 238726 88420
rect 289814 88408 289820 88420
rect 289872 88408 289878 88460
rect 293862 88408 293868 88460
rect 293920 88448 293926 88460
rect 345014 88448 345020 88460
rect 293920 88420 345020 88448
rect 293920 88408 293926 88420
rect 345014 88408 345020 88420
rect 345072 88408 345078 88460
rect 350442 88408 350448 88460
rect 350500 88448 350506 88460
rect 401594 88448 401600 88460
rect 350500 88420 401600 88448
rect 350500 88408 350506 88420
rect 401594 88408 401600 88420
rect 401652 88408 401658 88460
rect 434622 88408 434628 88460
rect 434680 88448 434686 88460
rect 485774 88448 485780 88460
rect 434680 88420 485780 88448
rect 434680 88408 434686 88420
rect 485774 88408 485780 88420
rect 485832 88408 485838 88460
rect 13722 88340 13728 88392
rect 13780 88380 13786 88392
rect 66254 88380 66260 88392
rect 13780 88352 66260 88380
rect 13780 88340 13786 88352
rect 66254 88340 66260 88352
rect 66312 88340 66318 88392
rect 70302 88340 70308 88392
rect 70360 88380 70366 88392
rect 121454 88380 121460 88392
rect 70360 88352 121460 88380
rect 70360 88340 70366 88352
rect 121454 88340 121460 88352
rect 121512 88340 121518 88392
rect 126882 88340 126888 88392
rect 126940 88380 126946 88392
rect 178034 88380 178040 88392
rect 126940 88352 178040 88380
rect 126940 88340 126946 88352
rect 178034 88340 178040 88352
rect 178092 88340 178098 88392
rect 209682 88340 209688 88392
rect 209740 88380 209746 88392
rect 262214 88380 262220 88392
rect 209740 88352 262220 88380
rect 209740 88340 209746 88352
rect 262214 88340 262220 88352
rect 262272 88340 262278 88392
rect 322842 88340 322848 88392
rect 322900 88380 322906 88392
rect 373994 88380 374000 88392
rect 322900 88352 374000 88380
rect 322900 88340 322906 88352
rect 373994 88340 374000 88352
rect 374052 88340 374058 88392
rect 405642 88340 405648 88392
rect 405700 88380 405706 88392
rect 458174 88380 458180 88392
rect 405700 88352 458180 88380
rect 405700 88340 405706 88352
rect 458174 88340 458180 88352
rect 458232 88340 458238 88392
rect 518802 88340 518808 88392
rect 518860 88380 518866 88392
rect 569954 88380 569960 88392
rect 518860 88352 569960 88380
rect 518860 88340 518866 88352
rect 569954 88340 569960 88352
rect 570012 88340 570018 88392
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 11790 84232 11796 84244
rect 3200 84204 11796 84232
rect 3200 84192 3206 84204
rect 11790 84192 11796 84204
rect 11848 84192 11854 84244
rect 428642 72428 428648 72480
rect 428700 72468 428706 72480
rect 435726 72468 435732 72480
rect 428700 72440 435732 72468
rect 428700 72428 428706 72440
rect 435726 72428 435732 72440
rect 435784 72428 435790 72480
rect 63586 72292 63592 72344
rect 63644 72332 63650 72344
rect 64322 72332 64328 72344
rect 63644 72304 64328 72332
rect 63644 72292 63650 72304
rect 64322 72292 64328 72304
rect 64380 72292 64386 72344
rect 232682 72292 232688 72344
rect 232740 72332 232746 72344
rect 239766 72332 239772 72344
rect 232740 72304 239772 72332
rect 232740 72292 232746 72304
rect 239766 72292 239772 72304
rect 239824 72292 239830 72344
rect 259730 72292 259736 72344
rect 259788 72332 259794 72344
rect 260190 72332 260196 72344
rect 259788 72304 260196 72332
rect 259788 72292 259794 72304
rect 260190 72292 260196 72304
rect 260248 72292 260254 72344
rect 316770 72292 316776 72344
rect 316828 72332 316834 72344
rect 323670 72332 323676 72344
rect 316828 72304 323676 72332
rect 316828 72292 316834 72304
rect 323670 72292 323676 72304
rect 323728 72292 323734 72344
rect 455690 72292 455696 72344
rect 455748 72332 455754 72344
rect 456150 72332 456156 72344
rect 455748 72304 456156 72332
rect 455748 72292 455754 72304
rect 456150 72292 456156 72304
rect 456208 72292 456214 72344
rect 483658 72224 483664 72276
rect 483716 72264 483722 72276
rect 491662 72264 491668 72276
rect 483716 72236 491668 72264
rect 483716 72224 483722 72236
rect 491662 72224 491668 72236
rect 491720 72224 491726 72276
rect 287698 72088 287704 72140
rect 287756 72128 287762 72140
rect 295702 72128 295708 72140
rect 287756 72100 295708 72128
rect 287756 72088 287762 72100
rect 295702 72088 295708 72100
rect 295760 72088 295766 72140
rect 512730 72088 512736 72140
rect 512788 72128 512794 72140
rect 519630 72128 519636 72140
rect 512788 72100 519636 72128
rect 512788 72088 512794 72100
rect 519630 72088 519636 72100
rect 519688 72088 519694 72140
rect 35618 71680 35624 71732
rect 35676 71720 35682 71732
rect 36906 71720 36912 71732
rect 35676 71692 36912 71720
rect 35676 71680 35682 71692
rect 36906 71680 36912 71692
rect 36964 71680 36970 71732
rect 97902 71680 97908 71732
rect 97960 71720 97966 71732
rect 149054 71720 149060 71732
rect 97960 71692 149060 71720
rect 97960 71680 97966 71692
rect 149054 71680 149060 71692
rect 149112 71680 149118 71732
rect 182082 71680 182088 71732
rect 182140 71720 182146 71732
rect 233234 71720 233240 71732
rect 182140 71692 233240 71720
rect 182140 71680 182146 71692
rect 233234 71680 233240 71692
rect 233292 71680 233298 71732
rect 266262 71680 266268 71732
rect 266320 71720 266326 71732
rect 317414 71720 317420 71732
rect 266320 71692 317420 71720
rect 266320 71680 266326 71692
rect 317414 71680 317420 71692
rect 317472 71680 317478 71732
rect 343542 71680 343548 71732
rect 343600 71720 343606 71732
rect 345658 71720 345664 71732
rect 343600 71692 345664 71720
rect 343600 71680 343606 71692
rect 345658 71680 345664 71692
rect 345716 71680 345722 71732
rect 378042 71680 378048 71732
rect 378100 71720 378106 71732
rect 429194 71720 429200 71732
rect 378100 71692 429200 71720
rect 378100 71680 378106 71692
rect 429194 71680 429200 71692
rect 429252 71680 429258 71732
rect 489822 71680 489828 71732
rect 489880 71720 489886 71732
rect 542354 71720 542360 71732
rect 489880 71692 542360 71720
rect 489880 71680 489886 71692
rect 542354 71680 542360 71692
rect 542412 71680 542418 71732
rect 231670 71612 231676 71664
rect 231728 71652 231734 71664
rect 232590 71652 232596 71664
rect 231728 71624 232596 71652
rect 231728 71612 231734 71624
rect 232590 71612 232596 71624
rect 232648 71612 232654 71664
rect 462222 71612 462228 71664
rect 462280 71652 462286 71664
rect 513374 71652 513380 71664
rect 462280 71624 513380 71652
rect 462280 71612 462286 71624
rect 513374 71612 513380 71624
rect 513432 71612 513438 71664
rect 42886 68960 42892 69012
rect 42944 69000 42950 69012
rect 72050 69000 72056 69012
rect 42944 68972 45554 69000
rect 42944 68960 42950 68972
rect 15194 68892 15200 68944
rect 15252 68932 15258 68944
rect 43990 68932 43996 68944
rect 15252 68904 43996 68932
rect 15252 68892 15258 68904
rect 43990 68892 43996 68904
rect 44048 68892 44054 68944
rect 45526 68932 45554 68972
rect 64846 68972 72056 69000
rect 64846 68932 64874 68972
rect 72050 68960 72056 68972
rect 72108 68960 72114 69012
rect 99466 68960 99472 69012
rect 99524 69000 99530 69012
rect 99524 68972 103514 69000
rect 99524 68960 99530 68972
rect 45526 68904 64874 68932
rect 71866 68892 71872 68944
rect 71924 68932 71930 68944
rect 100018 68932 100024 68944
rect 71924 68904 100024 68932
rect 71924 68892 71930 68904
rect 100018 68892 100024 68904
rect 100076 68892 100082 68944
rect 103486 68932 103514 68972
rect 127066 68960 127072 69012
rect 127124 69000 127130 69012
rect 127124 68972 132494 69000
rect 127124 68960 127130 68972
rect 127986 68932 127992 68944
rect 103486 68904 127992 68932
rect 127986 68892 127992 68904
rect 128044 68892 128050 68944
rect 132466 68932 132494 68972
rect 183646 68960 183652 69012
rect 183704 69000 183710 69012
rect 183704 68972 190454 69000
rect 183704 68960 183710 68972
rect 156046 68932 156052 68944
rect 132466 68904 156052 68932
rect 156046 68892 156052 68904
rect 156104 68892 156110 68944
rect 165982 68892 165988 68944
rect 166040 68932 166046 68944
rect 177298 68932 177304 68944
rect 166040 68904 177304 68932
rect 166040 68892 166046 68904
rect 177298 68892 177304 68904
rect 177356 68892 177362 68944
rect 178678 68892 178684 68944
rect 178736 68932 178742 68944
rect 184014 68932 184020 68944
rect 178736 68904 184020 68932
rect 178736 68892 178742 68904
rect 184014 68892 184020 68904
rect 184072 68892 184078 68944
rect 190426 68932 190454 68972
rect 374638 68960 374644 69012
rect 374696 69000 374702 69012
rect 379698 69000 379704 69012
rect 374696 68972 379704 69000
rect 374696 68960 374702 68972
rect 379698 68960 379704 68972
rect 379756 68960 379762 69012
rect 539318 68960 539324 69012
rect 539376 69000 539382 69012
rect 542998 69000 543004 69012
rect 539376 68972 543004 69000
rect 539376 68960 539382 68972
rect 542998 68960 543004 68972
rect 543056 68960 543062 69012
rect 211706 68932 211712 68944
rect 190426 68904 211712 68932
rect 211706 68892 211712 68904
rect 211764 68892 211770 68944
rect 222010 68892 222016 68944
rect 222068 68932 222074 68944
rect 232498 68932 232504 68944
rect 222068 68904 232504 68932
rect 222068 68892 222074 68904
rect 232498 68892 232504 68904
rect 232556 68892 232562 68944
rect 249702 68892 249708 68944
rect 249760 68932 249766 68944
rect 260098 68932 260104 68944
rect 249760 68904 260104 68932
rect 249760 68892 249766 68904
rect 260098 68892 260104 68904
rect 260156 68892 260162 68944
rect 261478 68892 261484 68944
rect 261536 68932 261542 68944
rect 567194 68932 567200 68944
rect 261536 68904 567200 68932
rect 261536 68892 261542 68904
rect 567194 68892 567200 68904
rect 567252 68892 567258 68944
rect 25682 68824 25688 68876
rect 25740 68864 25746 68876
rect 36998 68864 37004 68876
rect 25740 68836 37004 68864
rect 25740 68824 25746 68836
rect 36998 68824 37004 68836
rect 37056 68824 37062 68876
rect 53650 68824 53656 68876
rect 53708 68864 53714 68876
rect 69658 68864 69664 68876
rect 53708 68836 69664 68864
rect 53708 68824 53714 68836
rect 69658 68824 69664 68836
rect 69716 68824 69722 68876
rect 81986 68824 81992 68876
rect 82044 68864 82050 68876
rect 94498 68864 94504 68876
rect 82044 68836 94504 68864
rect 82044 68824 82050 68836
rect 94498 68824 94504 68836
rect 94556 68824 94562 68876
rect 109678 68824 109684 68876
rect 109736 68864 109742 68876
rect 120718 68864 120724 68876
rect 109736 68836 120724 68864
rect 109736 68824 109742 68836
rect 120718 68824 120724 68836
rect 120776 68824 120782 68876
rect 137646 68824 137652 68876
rect 137704 68864 137710 68876
rect 148410 68864 148416 68876
rect 137704 68836 148416 68864
rect 137704 68824 137710 68836
rect 148410 68824 148416 68836
rect 148468 68824 148474 68876
rect 193674 68824 193680 68876
rect 193732 68864 193738 68876
rect 204898 68864 204904 68876
rect 193732 68836 204904 68864
rect 193732 68824 193738 68836
rect 204898 68824 204904 68836
rect 204956 68824 204962 68876
rect 238846 68824 238852 68876
rect 238904 68864 238910 68876
rect 268010 68864 268016 68876
rect 238904 68836 268016 68864
rect 238904 68824 238910 68836
rect 268010 68824 268016 68836
rect 268068 68824 268074 68876
rect 277670 68824 277676 68876
rect 277728 68864 277734 68876
rect 289078 68864 289084 68876
rect 277728 68836 289084 68864
rect 277728 68824 277734 68836
rect 289078 68824 289084 68836
rect 289136 68824 289142 68876
rect 306006 68824 306012 68876
rect 306064 68864 306070 68876
rect 316678 68864 316684 68876
rect 306064 68836 316684 68864
rect 306064 68824 306070 68836
rect 316678 68824 316684 68836
rect 316736 68824 316742 68876
rect 323026 68824 323032 68876
rect 323084 68864 323090 68876
rect 352006 68864 352012 68876
rect 323084 68836 352012 68864
rect 323084 68824 323090 68836
rect 352006 68824 352012 68836
rect 352064 68824 352070 68876
rect 361666 68824 361672 68876
rect 361724 68864 361730 68876
rect 373258 68864 373264 68876
rect 361724 68836 373264 68864
rect 361724 68824 361730 68836
rect 373258 68824 373264 68836
rect 373316 68824 373322 68876
rect 379606 68824 379612 68876
rect 379664 68864 379670 68876
rect 408034 68864 408040 68876
rect 379664 68836 408040 68864
rect 379664 68824 379670 68836
rect 408034 68824 408040 68836
rect 408092 68824 408098 68876
rect 417694 68824 417700 68876
rect 417752 68864 417758 68876
rect 428550 68864 428556 68876
rect 417752 68836 428556 68864
rect 417752 68824 417758 68836
rect 428550 68824 428556 68836
rect 428608 68824 428614 68876
rect 434806 68824 434812 68876
rect 434864 68864 434870 68876
rect 463694 68864 463700 68876
rect 434864 68836 463700 68864
rect 434864 68824 434870 68836
rect 463694 68824 463700 68836
rect 463752 68824 463758 68876
rect 473998 68824 474004 68876
rect 474056 68864 474062 68876
rect 485038 68864 485044 68876
rect 474056 68836 485044 68864
rect 474056 68824 474062 68836
rect 485038 68824 485044 68836
rect 485096 68824 485102 68876
rect 501690 68824 501696 68876
rect 501748 68864 501754 68876
rect 512638 68864 512644 68876
rect 501748 68836 512644 68864
rect 501748 68824 501754 68836
rect 512638 68824 512644 68836
rect 512696 68824 512702 68876
rect 518986 68824 518992 68876
rect 519044 68864 519050 68876
rect 547874 68864 547880 68876
rect 519044 68836 547880 68864
rect 519044 68824 519050 68836
rect 547874 68824 547880 68836
rect 547932 68824 547938 68876
rect 333698 68756 333704 68808
rect 333756 68796 333762 68808
rect 344278 68796 344284 68808
rect 333756 68768 344284 68796
rect 333756 68756 333762 68768
rect 344278 68756 344284 68768
rect 344336 68756 344342 68808
rect 390002 68756 390008 68808
rect 390060 68796 390066 68808
rect 400858 68796 400864 68808
rect 390060 68768 400864 68796
rect 390060 68756 390066 68768
rect 400858 68756 400864 68768
rect 400916 68756 400922 68808
rect 445662 68756 445668 68808
rect 445720 68796 445726 68808
rect 456058 68796 456064 68808
rect 445720 68768 456064 68796
rect 445720 68756 445726 68768
rect 456058 68756 456064 68768
rect 456116 68756 456122 68808
rect 529658 68756 529664 68808
rect 529716 68796 529722 68808
rect 540238 68796 540244 68808
rect 529716 68768 540244 68796
rect 529716 68756 529722 68768
rect 540238 68756 540244 68768
rect 540296 68756 540302 68808
rect 36814 68688 36820 68740
rect 36872 68728 36878 68740
rect 557534 68728 557540 68740
rect 36872 68700 557540 68728
rect 36872 68688 36878 68700
rect 557534 68688 557540 68700
rect 557592 68688 557598 68740
rect 16022 65492 16028 65544
rect 16080 65532 16086 65544
rect 547874 65532 547880 65544
rect 16080 65504 547880 65532
rect 16080 65492 16086 65504
rect 547874 65492 547880 65504
rect 547932 65492 547938 65544
rect 25682 65152 25688 65204
rect 25740 65192 25746 65204
rect 261478 65192 261484 65204
rect 25740 65164 261484 65192
rect 25740 65152 25746 65164
rect 261478 65152 261484 65164
rect 261536 65152 261542 65204
rect 36906 65084 36912 65136
rect 36964 65124 36970 65136
rect 53650 65124 53656 65136
rect 36964 65096 53656 65124
rect 36964 65084 36970 65096
rect 53650 65084 53656 65096
rect 53708 65084 53714 65136
rect 148410 65084 148416 65136
rect 148468 65124 148474 65136
rect 165614 65124 165620 65136
rect 148468 65096 165620 65124
rect 148468 65084 148474 65096
rect 165614 65084 165620 65096
rect 165672 65084 165678 65136
rect 175458 65084 175464 65136
rect 175516 65124 175522 65136
rect 193674 65124 193680 65136
rect 175516 65096 193680 65124
rect 175516 65084 175522 65096
rect 193674 65084 193680 65096
rect 193732 65084 193738 65136
rect 203518 65084 203524 65136
rect 203576 65124 203582 65136
rect 221366 65124 221372 65136
rect 203576 65096 221372 65124
rect 203576 65084 203582 65096
rect 221366 65084 221372 65096
rect 221424 65084 221430 65136
rect 408034 65084 408040 65136
rect 408092 65124 408098 65136
rect 428642 65124 428648 65136
rect 408092 65096 428648 65124
rect 408092 65084 408098 65096
rect 428642 65084 428648 65096
rect 428700 65084 428706 65136
rect 36814 65016 36820 65068
rect 36872 65056 36878 65068
rect 63310 65056 63316 65068
rect 36872 65028 63316 65056
rect 36872 65016 36878 65028
rect 63310 65016 63316 65028
rect 63368 65016 63374 65068
rect 64414 65016 64420 65068
rect 64472 65056 64478 65068
rect 81434 65056 81440 65068
rect 64472 65028 81440 65056
rect 64472 65016 64478 65028
rect 81434 65016 81440 65028
rect 81492 65016 81498 65068
rect 91462 65016 91468 65068
rect 91520 65056 91526 65068
rect 109678 65056 109684 65068
rect 91520 65028 109684 65056
rect 91520 65016 91526 65028
rect 109678 65016 109684 65028
rect 109736 65016 109742 65068
rect 119430 65016 119436 65068
rect 119488 65056 119494 65068
rect 137646 65056 137652 65068
rect 119488 65028 137652 65056
rect 119488 65016 119494 65028
rect 137646 65016 137652 65028
rect 137704 65016 137710 65068
rect 156322 65016 156328 65068
rect 156380 65056 156386 65068
rect 178678 65056 178684 65068
rect 156380 65028 178684 65056
rect 156380 65016 156386 65028
rect 178678 65016 178684 65028
rect 178736 65016 178742 65068
rect 232498 65016 232504 65068
rect 232556 65056 232562 65068
rect 249702 65056 249708 65068
rect 232556 65028 249708 65056
rect 232556 65016 232562 65028
rect 249702 65016 249708 65028
rect 249760 65016 249766 65068
rect 260098 65016 260104 65068
rect 260156 65056 260162 65068
rect 277670 65056 277676 65068
rect 260156 65028 277676 65056
rect 260156 65016 260162 65028
rect 277670 65016 277676 65028
rect 277728 65016 277734 65068
rect 287514 65016 287520 65068
rect 287572 65056 287578 65068
rect 305362 65056 305368 65068
rect 287572 65028 305368 65056
rect 287572 65016 287578 65028
rect 305362 65016 305368 65028
rect 305420 65016 305426 65068
rect 315482 65016 315488 65068
rect 315540 65056 315546 65068
rect 333698 65056 333704 65068
rect 315540 65028 333704 65056
rect 315540 65016 315546 65028
rect 333698 65016 333704 65028
rect 333756 65016 333762 65068
rect 345658 65016 345664 65068
rect 345716 65056 345722 65068
rect 361666 65056 361672 65068
rect 345716 65028 361672 65056
rect 345716 65016 345722 65028
rect 361666 65016 361672 65028
rect 361724 65016 361730 65068
rect 371510 65016 371516 65068
rect 371568 65056 371574 65068
rect 389358 65056 389364 65068
rect 371568 65028 389364 65056
rect 371568 65016 371574 65028
rect 389358 65016 389364 65028
rect 389416 65016 389422 65068
rect 399478 65016 399484 65068
rect 399536 65056 399542 65068
rect 417694 65056 417700 65068
rect 399536 65028 417700 65056
rect 399536 65016 399542 65028
rect 417694 65016 417700 65028
rect 417752 65016 417758 65068
rect 456150 65016 456156 65068
rect 456208 65056 456214 65068
rect 473538 65056 473544 65068
rect 456208 65028 473544 65056
rect 456208 65016 456214 65028
rect 473538 65016 473544 65028
rect 473596 65016 473602 65068
rect 483474 65016 483480 65068
rect 483532 65056 483538 65068
rect 501690 65056 501696 65068
rect 483532 65028 501696 65056
rect 483532 65016 483538 65028
rect 501690 65016 501696 65028
rect 501748 65016 501754 65068
rect 511442 65016 511448 65068
rect 511500 65056 511506 65068
rect 529658 65056 529664 65068
rect 511500 65028 529664 65056
rect 511500 65016 511506 65028
rect 529658 65016 529664 65028
rect 529716 65016 529722 65068
rect 35342 64948 35348 65000
rect 35400 64988 35406 65000
rect 64322 64988 64328 65000
rect 35400 64960 64328 64988
rect 35400 64948 35406 64960
rect 64322 64948 64328 64960
rect 64380 64948 64386 65000
rect 66898 64948 66904 65000
rect 66956 64988 66962 65000
rect 91094 64988 91100 65000
rect 66956 64960 91100 64988
rect 66956 64948 66962 64960
rect 91094 64948 91100 64960
rect 91152 64948 91158 65000
rect 94498 64948 94504 65000
rect 94556 64988 94562 65000
rect 119338 64988 119344 65000
rect 94556 64960 119344 64988
rect 94556 64948 94562 64960
rect 119338 64948 119344 64960
rect 119396 64948 119402 65000
rect 120718 64948 120724 65000
rect 120776 64988 120782 65000
rect 147306 64988 147312 65000
rect 120776 64960 147312 64988
rect 120776 64948 120782 64960
rect 147306 64948 147312 64960
rect 147364 64948 147370 65000
rect 148318 64948 148324 65000
rect 148376 64988 148382 65000
rect 175274 64988 175280 65000
rect 148376 64960 175280 64988
rect 148376 64948 148382 64960
rect 175274 64948 175280 64960
rect 175332 64948 175338 65000
rect 177298 64948 177304 65000
rect 177356 64988 177362 65000
rect 203334 64988 203340 65000
rect 177356 64960 203340 64988
rect 177356 64948 177362 64960
rect 203334 64948 203340 64960
rect 203392 64948 203398 65000
rect 204898 64948 204904 65000
rect 204956 64988 204962 65000
rect 231026 64988 231032 65000
rect 204956 64960 231032 64988
rect 204956 64948 204962 64960
rect 231026 64948 231032 64960
rect 231084 64948 231090 65000
rect 232590 64948 232596 65000
rect 232648 64988 232654 65000
rect 259362 64988 259368 65000
rect 232648 64960 259368 64988
rect 232648 64948 232654 64960
rect 259362 64948 259368 64960
rect 259420 64948 259426 65000
rect 268010 64948 268016 65000
rect 268068 64988 268074 65000
rect 287698 64988 287704 65000
rect 268068 64960 287704 64988
rect 268068 64948 268074 64960
rect 287698 64948 287704 64960
rect 287756 64948 287762 65000
rect 296346 64948 296352 65000
rect 296404 64988 296410 65000
rect 316770 64988 316776 65000
rect 296404 64960 316776 64988
rect 296404 64948 296410 64960
rect 316770 64948 316776 64960
rect 316828 64948 316834 65000
rect 352006 64948 352012 65000
rect 352064 64988 352070 65000
rect 374638 64988 374644 65000
rect 352064 64960 374644 64988
rect 352064 64948 352070 64960
rect 374638 64948 374644 64960
rect 374696 64948 374702 65000
rect 428458 64948 428464 65000
rect 428516 64988 428522 65000
rect 445662 64988 445668 65000
rect 428516 64960 445668 64988
rect 428516 64948 428522 64960
rect 445662 64948 445668 64960
rect 445720 64948 445726 65000
rect 464338 64948 464344 65000
rect 464396 64988 464402 65000
rect 483658 64988 483664 65000
rect 464396 64960 483664 64988
rect 464396 64948 464402 64960
rect 483658 64948 483664 64960
rect 483716 64948 483722 65000
rect 492030 64948 492036 65000
rect 492088 64988 492094 65000
rect 512730 64988 512736 65000
rect 492088 64960 512736 64988
rect 492088 64948 492094 64960
rect 512730 64948 512736 64960
rect 512788 64948 512794 65000
rect 542998 64948 543004 65000
rect 543056 64988 543062 65000
rect 557534 64988 557540 65000
rect 543056 64960 557540 64988
rect 543056 64948 543062 64960
rect 557534 64948 557540 64960
rect 557592 64948 557598 65000
rect 212258 64880 212264 64932
rect 212316 64920 212322 64932
rect 232682 64920 232688 64932
rect 212316 64892 232688 64920
rect 212316 64880 212322 64892
rect 232682 64880 232688 64892
rect 232740 64880 232746 64932
rect 260190 64880 260196 64932
rect 260248 64920 260254 64932
rect 287330 64920 287336 64932
rect 260248 64892 287336 64920
rect 260248 64880 260254 64892
rect 287330 64880 287336 64892
rect 287388 64880 287394 64932
rect 289078 64880 289084 64932
rect 289136 64920 289142 64932
rect 315022 64920 315028 64932
rect 289136 64892 315028 64920
rect 289136 64880 289142 64892
rect 315022 64880 315028 64892
rect 315080 64880 315086 64932
rect 316678 64880 316684 64932
rect 316736 64920 316742 64932
rect 343358 64920 343364 64932
rect 316736 64892 343364 64920
rect 316736 64880 316742 64892
rect 343358 64880 343364 64892
rect 343416 64880 343422 64932
rect 344278 64880 344284 64932
rect 344336 64920 344342 64932
rect 371326 64920 371332 64932
rect 344336 64892 371332 64920
rect 344336 64880 344342 64892
rect 371326 64880 371332 64892
rect 371384 64880 371390 64932
rect 373258 64880 373264 64932
rect 373316 64920 373322 64932
rect 399018 64920 399024 64932
rect 373316 64892 399024 64920
rect 373316 64880 373322 64892
rect 399018 64880 399024 64892
rect 399076 64880 399082 64932
rect 400858 64880 400864 64932
rect 400916 64920 400922 64932
rect 427354 64920 427360 64932
rect 400916 64892 427360 64920
rect 400916 64880 400922 64892
rect 427354 64880 427360 64892
rect 427412 64880 427418 64932
rect 428550 64880 428556 64932
rect 428608 64920 428614 64932
rect 455322 64920 455328 64932
rect 428608 64892 455328 64920
rect 428608 64880 428614 64892
rect 455322 64880 455328 64892
rect 455380 64880 455386 64932
rect 456058 64880 456064 64932
rect 456116 64920 456122 64932
rect 483198 64920 483204 64932
rect 456116 64892 483204 64920
rect 456116 64880 456122 64892
rect 483198 64880 483204 64892
rect 483256 64880 483262 64932
rect 485038 64880 485044 64932
rect 485096 64920 485102 64932
rect 511350 64920 511356 64932
rect 485096 64892 511356 64920
rect 485096 64880 485102 64892
rect 511350 64880 511356 64892
rect 511408 64880 511414 64932
rect 512638 64880 512644 64932
rect 512696 64920 512702 64932
rect 539318 64920 539324 64932
rect 512696 64892 539324 64920
rect 512696 64880 512702 64892
rect 539318 64880 539324 64892
rect 539376 64880 539382 64932
rect 540238 64880 540244 64932
rect 540296 64920 540302 64932
rect 567194 64920 567200 64932
rect 540296 64892 567200 64920
rect 540296 64880 540302 64892
rect 567194 64880 567200 64892
rect 567252 64880 567258 64932
rect 37918 62772 37924 62824
rect 37976 62812 37982 62824
rect 545758 62812 545764 62824
rect 37976 62784 545764 62812
rect 37976 62772 37982 62784
rect 545758 62772 545764 62784
rect 545816 62772 545822 62824
rect 182082 62160 182088 62212
rect 182140 62200 182146 62212
rect 233234 62200 233240 62212
rect 182140 62172 233240 62200
rect 182140 62160 182146 62172
rect 233234 62160 233240 62172
rect 233292 62160 233298 62212
rect 350442 62160 350448 62212
rect 350500 62200 350506 62212
rect 401594 62200 401600 62212
rect 350500 62172 401600 62200
rect 350500 62160 350506 62172
rect 401594 62160 401600 62172
rect 401652 62160 401658 62212
rect 42702 62092 42708 62144
rect 42760 62132 42766 62144
rect 93854 62132 93860 62144
rect 42760 62104 93860 62132
rect 42760 62092 42766 62104
rect 93854 62092 93860 62104
rect 93912 62092 93918 62144
rect 97902 62092 97908 62144
rect 97960 62132 97966 62144
rect 149054 62132 149060 62144
rect 97960 62104 149060 62132
rect 97960 62092 97966 62104
rect 149054 62092 149060 62104
rect 149112 62092 149118 62144
rect 154482 62092 154488 62144
rect 154540 62132 154546 62144
rect 205634 62132 205640 62144
rect 154540 62104 205640 62132
rect 154540 62092 154546 62104
rect 205634 62092 205640 62104
rect 205692 62092 205698 62144
rect 238662 62092 238668 62144
rect 238720 62132 238726 62144
rect 289814 62132 289820 62144
rect 238720 62104 289820 62132
rect 238720 62092 238726 62104
rect 289814 62092 289820 62104
rect 289872 62092 289878 62144
rect 293862 62092 293868 62144
rect 293920 62132 293926 62144
rect 345014 62132 345020 62144
rect 293920 62104 345020 62132
rect 293920 62092 293926 62104
rect 345014 62092 345020 62104
rect 345072 62092 345078 62144
rect 378042 62092 378048 62144
rect 378100 62132 378106 62144
rect 429194 62132 429200 62144
rect 378100 62104 429200 62132
rect 378100 62092 378106 62104
rect 429194 62092 429200 62104
rect 429252 62092 429258 62144
rect 434622 62092 434628 62144
rect 434680 62132 434686 62144
rect 485774 62132 485780 62144
rect 434680 62104 485780 62132
rect 434680 62092 434686 62104
rect 485774 62092 485780 62104
rect 485832 62092 485838 62144
rect 489822 62092 489828 62144
rect 489880 62132 489886 62144
rect 542354 62132 542360 62144
rect 489880 62104 542360 62132
rect 489880 62092 489886 62104
rect 542354 62092 542360 62104
rect 542412 62092 542418 62144
rect 63586 50328 63592 50380
rect 63644 50368 63650 50380
rect 64414 50368 64420 50380
rect 63644 50340 64420 50368
rect 63644 50328 63650 50340
rect 64414 50328 64420 50340
rect 64472 50328 64478 50380
rect 147674 50328 147680 50380
rect 147732 50368 147738 50380
rect 148410 50368 148416 50380
rect 147732 50340 148416 50368
rect 147732 50328 147738 50340
rect 148410 50328 148416 50340
rect 148468 50328 148474 50380
rect 455690 50328 455696 50380
rect 455748 50368 455754 50380
rect 456150 50368 456156 50380
rect 455748 50340 456156 50368
rect 455748 50328 455754 50340
rect 456150 50328 456156 50340
rect 456208 50328 456214 50380
rect 232682 44888 232688 44940
rect 232740 44928 232746 44940
rect 239766 44928 239772 44940
rect 232740 44900 239772 44928
rect 232740 44888 232746 44900
rect 239766 44888 239772 44900
rect 239824 44888 239830 44940
rect 428642 44820 428648 44872
rect 428700 44860 428706 44872
rect 435726 44860 435732 44872
rect 428700 44832 435732 44860
rect 428700 44820 428706 44832
rect 435726 44820 435732 44832
rect 435784 44820 435790 44872
rect 512730 44684 512736 44736
rect 512788 44724 512794 44736
rect 519630 44724 519636 44736
rect 512788 44696 519636 44724
rect 512788 44684 512794 44696
rect 519630 44684 519636 44696
rect 519688 44684 519694 44736
rect 483658 44616 483664 44668
rect 483716 44656 483722 44668
rect 491662 44656 491668 44668
rect 483716 44628 491668 44656
rect 483716 44616 483722 44628
rect 491662 44616 491668 44628
rect 491720 44616 491726 44668
rect 3234 44480 3240 44532
rect 3292 44520 3298 44532
rect 8938 44520 8944 44532
rect 3292 44492 8944 44520
rect 3292 44480 3298 44492
rect 8938 44480 8944 44492
rect 8996 44480 9002 44532
rect 287698 44276 287704 44328
rect 287756 44316 287762 44328
rect 295702 44316 295708 44328
rect 287756 44288 295708 44316
rect 287756 44276 287762 44288
rect 295702 44276 295708 44288
rect 295760 44276 295766 44328
rect 316770 44276 316776 44328
rect 316828 44316 316834 44328
rect 323670 44316 323676 44328
rect 316828 44288 323676 44316
rect 316828 44276 316834 44288
rect 323670 44276 323676 44288
rect 323728 44276 323734 44328
rect 13722 44072 13728 44124
rect 13780 44112 13786 44124
rect 66254 44112 66260 44124
rect 13780 44084 66260 44112
rect 13780 44072 13786 44084
rect 66254 44072 66260 44084
rect 66312 44072 66318 44124
rect 70302 44072 70308 44124
rect 70360 44112 70366 44124
rect 121454 44112 121460 44124
rect 70360 44084 121460 44112
rect 70360 44072 70366 44084
rect 121454 44072 121460 44084
rect 121512 44072 121518 44124
rect 126882 44072 126888 44124
rect 126940 44112 126946 44124
rect 178034 44112 178040 44124
rect 126940 44084 178040 44112
rect 126940 44072 126946 44084
rect 178034 44072 178040 44084
rect 178092 44072 178098 44124
rect 209682 44072 209688 44124
rect 209740 44112 209746 44124
rect 262214 44112 262220 44124
rect 209740 44084 262220 44112
rect 209740 44072 209746 44084
rect 262214 44072 262220 44084
rect 262272 44072 262278 44124
rect 266262 44072 266268 44124
rect 266320 44112 266326 44124
rect 317414 44112 317420 44124
rect 266320 44084 317420 44112
rect 266320 44072 266326 44084
rect 317414 44072 317420 44084
rect 317472 44072 317478 44124
rect 322842 44072 322848 44124
rect 322900 44112 322906 44124
rect 373994 44112 374000 44124
rect 322900 44084 374000 44112
rect 322900 44072 322906 44084
rect 373994 44072 374000 44084
rect 374052 44072 374058 44124
rect 405642 44072 405648 44124
rect 405700 44112 405706 44124
rect 458174 44112 458180 44124
rect 405700 44084 458180 44112
rect 405700 44072 405706 44084
rect 458174 44072 458180 44084
rect 458232 44072 458238 44124
rect 462222 44072 462228 44124
rect 462280 44112 462286 44124
rect 513374 44112 513380 44124
rect 462280 44084 513380 44112
rect 462280 44072 462286 44084
rect 513374 44072 513380 44084
rect 513432 44072 513438 44124
rect 518802 44072 518808 44124
rect 518860 44112 518866 44124
rect 569954 44112 569960 44124
rect 518860 44084 569960 44112
rect 518860 44072 518866 44084
rect 569954 44072 569960 44084
rect 570012 44072 570018 44124
rect 35618 44004 35624 44056
rect 35676 44044 35682 44056
rect 36906 44044 36912 44056
rect 35676 44016 36912 44044
rect 35676 44004 35682 44016
rect 36906 44004 36912 44016
rect 36964 44004 36970 44056
rect 343542 44004 343548 44056
rect 343600 44044 343606 44056
rect 345658 44044 345664 44056
rect 343600 44016 345664 44044
rect 343600 44004 343606 44016
rect 345658 44004 345664 44016
rect 345716 44004 345722 44056
rect 539502 44004 539508 44056
rect 539560 44044 539566 44056
rect 542998 44044 543004 44056
rect 539560 44016 543004 44044
rect 539560 44004 539566 44016
rect 542998 44004 543004 44016
rect 543056 44004 543062 44056
rect 25682 41352 25688 41404
rect 25740 41392 25746 41404
rect 36814 41392 36820 41404
rect 25740 41364 36820 41392
rect 25740 41352 25746 41364
rect 36814 41352 36820 41364
rect 36872 41352 36878 41404
rect 178678 41352 178684 41404
rect 178736 41392 178742 41404
rect 184014 41392 184020 41404
rect 178736 41364 184020 41392
rect 178736 41352 178742 41364
rect 184014 41352 184020 41364
rect 184072 41352 184078 41404
rect 374638 41352 374644 41404
rect 374696 41392 374702 41404
rect 379698 41392 379704 41404
rect 374696 41364 379704 41392
rect 374696 41352 374702 41364
rect 379698 41352 379704 41364
rect 379756 41352 379762 41404
rect 15194 41284 15200 41336
rect 15252 41324 15258 41336
rect 43990 41324 43996 41336
rect 15252 41296 43996 41324
rect 15252 41284 15258 41296
rect 43990 41284 43996 41296
rect 44048 41284 44054 41336
rect 71038 41284 71044 41336
rect 71096 41324 71102 41336
rect 567194 41324 567200 41336
rect 71096 41296 567200 41324
rect 71096 41284 71102 41296
rect 567194 41284 567200 41296
rect 567252 41284 567258 41336
rect 53650 41216 53656 41268
rect 53708 41256 53714 41268
rect 66898 41256 66904 41268
rect 53708 41228 66904 41256
rect 53708 41216 53714 41228
rect 66898 41216 66904 41228
rect 66956 41216 66962 41268
rect 71866 41216 71872 41268
rect 71924 41256 71930 41268
rect 100018 41256 100024 41268
rect 71924 41228 100024 41256
rect 71924 41216 71930 41228
rect 100018 41216 100024 41228
rect 100076 41216 100082 41268
rect 127986 41256 127992 41268
rect 103486 41228 127992 41256
rect 42886 41148 42892 41200
rect 42944 41188 42950 41200
rect 72050 41188 72056 41200
rect 42944 41160 72056 41188
rect 42944 41148 42950 41160
rect 72050 41148 72056 41160
rect 72108 41148 72114 41200
rect 81986 41148 81992 41200
rect 82044 41188 82050 41200
rect 94498 41188 94504 41200
rect 82044 41160 94504 41188
rect 82044 41148 82050 41160
rect 94498 41148 94504 41160
rect 94556 41148 94562 41200
rect 99466 41148 99472 41200
rect 99524 41188 99530 41200
rect 103486 41188 103514 41228
rect 127986 41216 127992 41228
rect 128044 41216 128050 41268
rect 156046 41256 156052 41268
rect 132466 41228 156052 41256
rect 99524 41160 103514 41188
rect 99524 41148 99530 41160
rect 109678 41148 109684 41200
rect 109736 41188 109742 41200
rect 120718 41188 120724 41200
rect 109736 41160 120724 41188
rect 109736 41148 109742 41160
rect 120718 41148 120724 41160
rect 120776 41148 120782 41200
rect 127066 41148 127072 41200
rect 127124 41188 127130 41200
rect 132466 41188 132494 41228
rect 156046 41216 156052 41228
rect 156104 41216 156110 41268
rect 165982 41216 165988 41268
rect 166040 41256 166046 41268
rect 177298 41256 177304 41268
rect 166040 41228 177304 41256
rect 166040 41216 166046 41228
rect 177298 41216 177304 41228
rect 177356 41216 177362 41268
rect 183646 41216 183652 41268
rect 183704 41256 183710 41268
rect 211706 41256 211712 41268
rect 183704 41228 211712 41256
rect 183704 41216 183710 41228
rect 211706 41216 211712 41228
rect 211764 41216 211770 41268
rect 222010 41216 222016 41268
rect 222068 41256 222074 41268
rect 232590 41256 232596 41268
rect 222068 41228 232596 41256
rect 222068 41216 222074 41228
rect 232590 41216 232596 41228
rect 232648 41216 232654 41268
rect 238846 41216 238852 41268
rect 238904 41256 238910 41268
rect 268010 41256 268016 41268
rect 238904 41228 268016 41256
rect 238904 41216 238910 41228
rect 268010 41216 268016 41228
rect 268068 41216 268074 41268
rect 277670 41216 277676 41268
rect 277728 41256 277734 41268
rect 289078 41256 289084 41268
rect 277728 41228 289084 41256
rect 277728 41216 277734 41228
rect 289078 41216 289084 41228
rect 289136 41216 289142 41268
rect 306006 41216 306012 41268
rect 306064 41256 306070 41268
rect 316678 41256 316684 41268
rect 306064 41228 316684 41256
rect 306064 41216 306070 41228
rect 316678 41216 316684 41228
rect 316736 41216 316742 41268
rect 323026 41216 323032 41268
rect 323084 41256 323090 41268
rect 352006 41256 352012 41268
rect 323084 41228 352012 41256
rect 323084 41216 323090 41228
rect 352006 41216 352012 41228
rect 352064 41216 352070 41268
rect 361666 41216 361672 41268
rect 361724 41256 361730 41268
rect 373258 41256 373264 41268
rect 361724 41228 373264 41256
rect 361724 41216 361730 41228
rect 373258 41216 373264 41228
rect 373316 41216 373322 41268
rect 379606 41216 379612 41268
rect 379664 41256 379670 41268
rect 408034 41256 408040 41268
rect 379664 41228 408040 41256
rect 379664 41216 379670 41228
rect 408034 41216 408040 41228
rect 408092 41216 408098 41268
rect 417694 41216 417700 41268
rect 417752 41256 417758 41268
rect 428550 41256 428556 41268
rect 417752 41228 428556 41256
rect 417752 41216 417758 41228
rect 428550 41216 428556 41228
rect 428608 41216 428614 41268
rect 434806 41216 434812 41268
rect 434864 41256 434870 41268
rect 463694 41256 463700 41268
rect 434864 41228 463700 41256
rect 434864 41216 434870 41228
rect 463694 41216 463700 41228
rect 463752 41216 463758 41268
rect 473998 41216 474004 41268
rect 474056 41256 474062 41268
rect 485038 41256 485044 41268
rect 474056 41228 485044 41256
rect 474056 41216 474062 41228
rect 485038 41216 485044 41228
rect 485096 41216 485102 41268
rect 501690 41216 501696 41268
rect 501748 41256 501754 41268
rect 512638 41256 512644 41268
rect 501748 41228 512644 41256
rect 501748 41216 501754 41228
rect 512638 41216 512644 41228
rect 512696 41216 512702 41268
rect 518986 41216 518992 41268
rect 519044 41256 519050 41268
rect 547874 41256 547880 41268
rect 519044 41228 547880 41256
rect 519044 41216 519050 41228
rect 547874 41216 547880 41228
rect 547932 41216 547938 41268
rect 127124 41160 132494 41188
rect 127124 41148 127130 41160
rect 137646 41148 137652 41200
rect 137704 41188 137710 41200
rect 148318 41188 148324 41200
rect 137704 41160 148324 41188
rect 137704 41148 137710 41160
rect 148318 41148 148324 41160
rect 148376 41148 148382 41200
rect 193674 41148 193680 41200
rect 193732 41188 193738 41200
rect 204898 41188 204904 41200
rect 193732 41160 204904 41188
rect 193732 41148 193738 41160
rect 204898 41148 204904 41160
rect 204956 41148 204962 41200
rect 249702 41148 249708 41200
rect 249760 41188 249766 41200
rect 260190 41188 260196 41200
rect 249760 41160 260196 41188
rect 249760 41148 249766 41160
rect 260190 41148 260196 41160
rect 260248 41148 260254 41200
rect 333698 41148 333704 41200
rect 333756 41188 333762 41200
rect 344278 41188 344284 41200
rect 333756 41160 344284 41188
rect 333756 41148 333762 41160
rect 344278 41148 344284 41160
rect 344336 41148 344342 41200
rect 390002 41148 390008 41200
rect 390060 41188 390066 41200
rect 400858 41188 400864 41200
rect 390060 41160 400864 41188
rect 390060 41148 390066 41160
rect 400858 41148 400864 41160
rect 400916 41148 400922 41200
rect 445662 41148 445668 41200
rect 445720 41188 445726 41200
rect 456058 41188 456064 41200
rect 445720 41160 456064 41188
rect 445720 41148 445726 41160
rect 456058 41148 456064 41160
rect 456116 41148 456122 41200
rect 529658 41148 529664 41200
rect 529716 41188 529722 41200
rect 540238 41188 540244 41200
rect 529716 41160 540244 41188
rect 529716 41148 529722 41160
rect 540238 41148 540244 41160
rect 540296 41148 540302 41200
rect 36722 41080 36728 41132
rect 36780 41120 36786 41132
rect 557534 41120 557540 41132
rect 36780 41092 557540 41120
rect 36780 41080 36786 41092
rect 557534 41080 557540 41092
rect 557592 41080 557598 41132
rect 21174 38360 21180 38412
rect 21232 38400 21238 38412
rect 36538 38400 36544 38412
rect 21232 38372 36544 38400
rect 21232 38360 21238 38372
rect 36538 38360 36544 38372
rect 36596 38360 36602 38412
rect 11790 38292 11796 38344
rect 11848 38332 11854 38344
rect 34054 38332 34060 38344
rect 11848 38304 34060 38332
rect 11848 38292 11854 38304
rect 34054 38292 34060 38304
rect 34112 38292 34118 38344
rect 40034 38292 40040 38344
rect 40092 38332 40098 38344
rect 60734 38332 60740 38344
rect 40092 38304 60740 38332
rect 40092 38292 40098 38304
rect 60734 38292 60740 38304
rect 60792 38292 60798 38344
rect 13078 38224 13084 38276
rect 13136 38264 13142 38276
rect 52730 38264 52736 38276
rect 13136 38236 52736 38264
rect 13136 38224 13142 38236
rect 52730 38224 52736 38236
rect 52788 38224 52794 38276
rect 3418 38156 3424 38208
rect 3476 38196 3482 38208
rect 49510 38196 49516 38208
rect 3476 38168 49516 38196
rect 3476 38156 3482 38168
rect 49510 38156 49516 38168
rect 49568 38156 49574 38208
rect 3510 38088 3516 38140
rect 3568 38128 3574 38140
rect 59170 38128 59176 38140
rect 3568 38100 59176 38128
rect 3568 38088 3574 38100
rect 59170 38088 59176 38100
rect 59228 38088 59234 38140
rect 6178 38020 6184 38072
rect 6236 38060 6242 38072
rect 17954 38060 17960 38072
rect 6236 38032 17960 38060
rect 6236 38020 6242 38032
rect 17954 38020 17960 38032
rect 18012 38020 18018 38072
rect 24394 38020 24400 38072
rect 24452 38060 24458 38072
rect 234614 38060 234620 38072
rect 24452 38032 234620 38060
rect 24452 38020 24458 38032
rect 234614 38020 234620 38032
rect 234672 38020 234678 38072
rect 3694 37952 3700 38004
rect 3752 37992 3758 38004
rect 37274 37992 37280 38004
rect 3752 37964 37280 37992
rect 3752 37952 3758 37964
rect 37274 37952 37280 37964
rect 37332 37952 37338 38004
rect 46290 37952 46296 38004
rect 46348 37992 46354 38004
rect 567838 37992 567844 38004
rect 46348 37964 567844 37992
rect 46348 37952 46354 37964
rect 567838 37952 567844 37964
rect 567896 37952 567902 38004
rect 16022 37884 16028 37936
rect 16080 37924 16086 37936
rect 547966 37924 547972 37936
rect 16080 37896 547972 37924
rect 16080 37884 16086 37896
rect 547966 37884 547972 37896
rect 548024 37884 548030 37936
rect 212350 37476 212356 37528
rect 212408 37516 212414 37528
rect 232682 37516 232688 37528
rect 212408 37488 232688 37516
rect 212408 37476 212414 37488
rect 232682 37476 232688 37488
rect 232740 37476 232746 37528
rect 408034 37476 408040 37528
rect 408092 37516 408098 37528
rect 428642 37516 428648 37528
rect 408092 37488 428648 37516
rect 408092 37476 408098 37488
rect 428642 37476 428648 37488
rect 428700 37476 428706 37528
rect 30834 37408 30840 37460
rect 30892 37448 30898 37460
rect 36630 37448 36636 37460
rect 30892 37420 36636 37448
rect 30892 37408 30898 37420
rect 36630 37408 36636 37420
rect 36688 37408 36694 37460
rect 148318 37408 148324 37460
rect 148376 37448 148382 37460
rect 165706 37448 165712 37460
rect 148376 37420 165712 37448
rect 148376 37408 148382 37420
rect 165706 37408 165712 37420
rect 165764 37408 165770 37460
rect 175458 37408 175464 37460
rect 175516 37448 175522 37460
rect 193674 37448 193680 37460
rect 175516 37420 193680 37448
rect 175516 37408 175522 37420
rect 193674 37408 193680 37420
rect 193732 37408 193738 37460
rect 203518 37408 203524 37460
rect 203576 37448 203582 37460
rect 221366 37448 221372 37460
rect 203576 37420 221372 37448
rect 203576 37408 203582 37420
rect 221366 37408 221372 37420
rect 221424 37408 221430 37460
rect 260190 37408 260196 37460
rect 260248 37448 260254 37460
rect 277670 37448 277676 37460
rect 260248 37420 277676 37448
rect 260248 37408 260254 37420
rect 277670 37408 277676 37420
rect 277728 37408 277734 37460
rect 287514 37408 287520 37460
rect 287572 37448 287578 37460
rect 305362 37448 305368 37460
rect 287572 37420 305368 37448
rect 287572 37408 287578 37420
rect 305362 37408 305368 37420
rect 305420 37408 305426 37460
rect 345658 37408 345664 37460
rect 345716 37448 345722 37460
rect 361666 37448 361672 37460
rect 345716 37420 361672 37448
rect 345716 37408 345722 37420
rect 361666 37408 361672 37420
rect 361724 37408 361730 37460
rect 371510 37408 371516 37460
rect 371568 37448 371574 37460
rect 389358 37448 389364 37460
rect 371568 37420 389364 37448
rect 371568 37408 371574 37420
rect 389358 37408 389364 37420
rect 389416 37408 389422 37460
rect 399478 37408 399484 37460
rect 399536 37448 399542 37460
rect 417694 37448 417700 37460
rect 399536 37420 417700 37448
rect 399536 37408 399542 37420
rect 417694 37408 417700 37420
rect 417752 37408 417758 37460
rect 456058 37408 456064 37460
rect 456116 37448 456122 37460
rect 473354 37448 473360 37460
rect 456116 37420 473360 37448
rect 456116 37408 456122 37420
rect 473354 37408 473360 37420
rect 473412 37408 473418 37460
rect 483474 37408 483480 37460
rect 483532 37448 483538 37460
rect 501690 37448 501696 37460
rect 483532 37420 501696 37448
rect 483532 37408 483538 37420
rect 501690 37408 501696 37420
rect 501748 37408 501754 37460
rect 27614 37340 27620 37392
rect 27672 37380 27678 37392
rect 62758 37380 62764 37392
rect 27672 37352 62764 37380
rect 27672 37340 27678 37352
rect 62758 37340 62764 37352
rect 62816 37340 62822 37392
rect 64414 37340 64420 37392
rect 64472 37380 64478 37392
rect 81434 37380 81440 37392
rect 64472 37352 81440 37380
rect 64472 37340 64478 37352
rect 81434 37340 81440 37352
rect 81492 37340 81498 37392
rect 91462 37340 91468 37392
rect 91520 37380 91526 37392
rect 109678 37380 109684 37392
rect 91520 37352 109684 37380
rect 91520 37340 91526 37352
rect 109678 37340 109684 37352
rect 109736 37340 109742 37392
rect 126238 37340 126244 37392
rect 126296 37380 126302 37392
rect 137646 37380 137652 37392
rect 126296 37352 137652 37380
rect 126296 37340 126302 37352
rect 137646 37340 137652 37352
rect 137704 37340 137710 37392
rect 156322 37340 156328 37392
rect 156380 37380 156386 37392
rect 178678 37380 178684 37392
rect 156380 37352 178684 37380
rect 156380 37340 156386 37352
rect 178678 37340 178684 37352
rect 178736 37340 178742 37392
rect 232590 37340 232596 37392
rect 232648 37380 232654 37392
rect 249702 37380 249708 37392
rect 232648 37352 249708 37380
rect 232648 37340 232654 37352
rect 249702 37340 249708 37352
rect 249760 37340 249766 37392
rect 268010 37340 268016 37392
rect 268068 37380 268074 37392
rect 287698 37380 287704 37392
rect 268068 37352 287704 37380
rect 268068 37340 268074 37352
rect 287698 37340 287704 37352
rect 287756 37340 287762 37392
rect 296162 37340 296168 37392
rect 296220 37380 296226 37392
rect 316770 37380 316776 37392
rect 296220 37352 316776 37380
rect 296220 37340 296226 37352
rect 316770 37340 316776 37352
rect 316828 37340 316834 37392
rect 322198 37340 322204 37392
rect 322256 37380 322262 37392
rect 333698 37380 333704 37392
rect 322256 37352 333704 37380
rect 322256 37340 322262 37352
rect 333698 37340 333704 37352
rect 333756 37340 333762 37392
rect 352006 37340 352012 37392
rect 352064 37380 352070 37392
rect 374638 37380 374644 37392
rect 352064 37352 374644 37380
rect 352064 37340 352070 37352
rect 374638 37340 374644 37352
rect 374696 37340 374702 37392
rect 428458 37340 428464 37392
rect 428516 37380 428522 37392
rect 445662 37380 445668 37392
rect 428516 37352 445668 37380
rect 428516 37340 428522 37352
rect 445662 37340 445668 37352
rect 445720 37340 445726 37392
rect 464338 37340 464344 37392
rect 464396 37380 464402 37392
rect 483658 37380 483664 37392
rect 464396 37352 483664 37380
rect 464396 37340 464402 37352
rect 483658 37340 483664 37352
rect 483716 37340 483722 37392
rect 492030 37340 492036 37392
rect 492088 37380 492094 37392
rect 512730 37380 512736 37392
rect 492088 37352 512736 37380
rect 492088 37340 492094 37352
rect 512730 37340 512736 37352
rect 512788 37340 512794 37392
rect 518158 37340 518164 37392
rect 518216 37380 518222 37392
rect 529658 37380 529664 37392
rect 518216 37352 529664 37380
rect 518216 37340 518222 37352
rect 529658 37340 529664 37352
rect 529716 37340 529722 37392
rect 542998 37340 543004 37392
rect 543056 37380 543062 37392
rect 557534 37380 557540 37392
rect 543056 37352 557540 37380
rect 543056 37340 543062 37352
rect 557534 37340 557540 37352
rect 557592 37340 557598 37392
rect 1394 37272 1400 37324
rect 1452 37312 1458 37324
rect 39850 37312 39856 37324
rect 1452 37284 39856 37312
rect 1452 37272 1458 37284
rect 39850 37272 39856 37284
rect 39908 37272 39914 37324
rect 43070 37272 43076 37324
rect 43128 37312 43134 37324
rect 91094 37312 91100 37324
rect 43128 37284 91100 37312
rect 43128 37272 43134 37284
rect 91094 37272 91100 37284
rect 91152 37272 91158 37324
rect 93118 37272 93124 37324
rect 93176 37312 93182 37324
rect 119338 37312 119344 37324
rect 93176 37284 119344 37312
rect 93176 37272 93182 37284
rect 119338 37272 119344 37284
rect 119396 37272 119402 37324
rect 120718 37272 120724 37324
rect 120776 37312 120782 37324
rect 147306 37312 147312 37324
rect 120776 37284 147312 37312
rect 120776 37272 120782 37284
rect 147306 37272 147312 37284
rect 147364 37272 147370 37324
rect 148410 37272 148416 37324
rect 148468 37312 148474 37324
rect 175366 37312 175372 37324
rect 148468 37284 175372 37312
rect 148468 37272 148474 37284
rect 175366 37272 175372 37284
rect 175424 37272 175430 37324
rect 177298 37272 177304 37324
rect 177356 37312 177362 37324
rect 203334 37312 203340 37324
rect 177356 37284 203340 37312
rect 177356 37272 177362 37284
rect 203334 37272 203340 37284
rect 203392 37272 203398 37324
rect 204898 37272 204904 37324
rect 204956 37312 204962 37324
rect 231026 37312 231032 37324
rect 204956 37284 231032 37312
rect 204956 37272 204962 37284
rect 231026 37272 231032 37284
rect 231084 37272 231090 37324
rect 232498 37272 232504 37324
rect 232556 37312 232562 37324
rect 259362 37312 259368 37324
rect 232556 37284 259368 37312
rect 232556 37272 232562 37284
rect 259362 37272 259368 37284
rect 259420 37272 259426 37324
rect 260098 37272 260104 37324
rect 260156 37312 260162 37324
rect 287330 37312 287336 37324
rect 260156 37284 287336 37312
rect 260156 37272 260162 37284
rect 287330 37272 287336 37284
rect 287388 37272 287394 37324
rect 289078 37272 289084 37324
rect 289136 37312 289142 37324
rect 315022 37312 315028 37324
rect 289136 37284 315028 37312
rect 289136 37272 289142 37284
rect 315022 37272 315028 37284
rect 315080 37272 315086 37324
rect 316678 37272 316684 37324
rect 316736 37312 316742 37324
rect 343358 37312 343364 37324
rect 316736 37284 343364 37312
rect 316736 37272 316742 37284
rect 343358 37272 343364 37284
rect 343416 37272 343422 37324
rect 344278 37272 344284 37324
rect 344336 37312 344342 37324
rect 371326 37312 371332 37324
rect 344336 37284 371332 37312
rect 344336 37272 344342 37284
rect 371326 37272 371332 37284
rect 371384 37272 371390 37324
rect 373258 37272 373264 37324
rect 373316 37312 373322 37324
rect 399018 37312 399024 37324
rect 373316 37284 399024 37312
rect 373316 37272 373322 37284
rect 399018 37272 399024 37284
rect 399076 37272 399082 37324
rect 400858 37272 400864 37324
rect 400916 37312 400922 37324
rect 427354 37312 427360 37324
rect 400916 37284 427360 37312
rect 400916 37272 400922 37284
rect 427354 37272 427360 37284
rect 427412 37272 427418 37324
rect 428550 37272 428556 37324
rect 428608 37312 428614 37324
rect 455322 37312 455328 37324
rect 428608 37284 455328 37312
rect 428608 37272 428614 37284
rect 455322 37272 455328 37284
rect 455380 37272 455386 37324
rect 456150 37272 456156 37324
rect 456208 37312 456214 37324
rect 483014 37312 483020 37324
rect 456208 37284 483020 37312
rect 456208 37272 456214 37284
rect 483014 37272 483020 37284
rect 483072 37272 483078 37324
rect 485038 37272 485044 37324
rect 485096 37312 485102 37324
rect 511350 37312 511356 37324
rect 485096 37284 511356 37312
rect 485096 37272 485102 37284
rect 511350 37272 511356 37284
rect 511408 37272 511414 37324
rect 512638 37272 512644 37324
rect 512696 37312 512702 37324
rect 539318 37312 539324 37324
rect 512696 37284 539324 37312
rect 512696 37272 512702 37284
rect 539318 37272 539324 37284
rect 539376 37272 539382 37324
rect 547138 37272 547144 37324
rect 547196 37312 547202 37324
rect 567194 37312 567200 37324
rect 547196 37284 567200 37312
rect 547196 37272 547202 37284
rect 567194 37272 567200 37284
rect 567252 37272 567258 37324
rect 3970 36796 3976 36848
rect 4028 36836 4034 36848
rect 63678 36836 63684 36848
rect 4028 36808 63684 36836
rect 4028 36796 4034 36808
rect 63678 36796 63684 36808
rect 63736 36796 63742 36848
rect 3602 36728 3608 36780
rect 3660 36768 3666 36780
rect 63586 36768 63592 36780
rect 3660 36740 63592 36768
rect 3660 36728 3666 36740
rect 63586 36728 63592 36740
rect 63644 36728 63650 36780
rect 3326 36660 3332 36712
rect 3384 36700 3390 36712
rect 63494 36700 63500 36712
rect 3384 36672 63500 36700
rect 3384 36660 3390 36672
rect 63494 36660 63500 36672
rect 63552 36660 63558 36712
rect 37918 36592 37924 36644
rect 37976 36632 37982 36644
rect 545758 36632 545764 36644
rect 37976 36604 545764 36632
rect 37976 36592 37982 36604
rect 545758 36592 545764 36604
rect 545816 36592 545822 36644
rect 13630 36524 13636 36576
rect 13688 36564 13694 36576
rect 580258 36564 580264 36576
rect 13688 36536 580264 36564
rect 13688 36524 13694 36536
rect 580258 36524 580264 36536
rect 580316 36524 580322 36576
rect 3418 36048 3424 36100
rect 3476 36088 3482 36100
rect 61286 36088 61292 36100
rect 3476 36060 61292 36088
rect 3476 36048 3482 36060
rect 61286 36048 61292 36060
rect 61344 36048 61350 36100
rect 13722 35980 13728 36032
rect 13780 36020 13786 36032
rect 93854 36020 93860 36032
rect 13780 35992 93860 36020
rect 13780 35980 13786 35992
rect 93854 35980 93860 35992
rect 93912 35980 93918 36032
rect 14 35912 20 35964
rect 72 35952 78 35964
rect 55582 35952 55588 35964
rect 72 35924 55588 35952
rect 72 35912 78 35924
rect 55582 35912 55588 35924
rect 55640 35912 55646 35964
rect 126882 34620 126888 34672
rect 126940 34660 126946 34672
rect 178034 34660 178040 34672
rect 126940 34632 178040 34660
rect 126940 34620 126946 34632
rect 178034 34620 178040 34632
rect 178092 34620 178098 34672
rect 350442 34620 350448 34672
rect 350500 34660 350506 34672
rect 401594 34660 401600 34672
rect 350500 34632 401600 34660
rect 350500 34620 350506 34632
rect 401594 34620 401600 34632
rect 401652 34620 401658 34672
rect 434622 34620 434628 34672
rect 434680 34660 434686 34672
rect 485774 34660 485780 34672
rect 434680 34632 485780 34660
rect 434680 34620 434686 34632
rect 485774 34620 485780 34632
rect 485832 34620 485838 34672
rect 97902 34552 97908 34604
rect 97960 34592 97966 34604
rect 149054 34592 149060 34604
rect 97960 34564 149060 34592
rect 97960 34552 97966 34564
rect 149054 34552 149060 34564
rect 149112 34552 149118 34604
rect 182082 34552 182088 34604
rect 182140 34592 182146 34604
rect 233234 34592 233240 34604
rect 182140 34564 233240 34592
rect 182140 34552 182146 34564
rect 233234 34552 233240 34564
rect 233292 34552 233298 34604
rect 238662 34552 238668 34604
rect 238720 34592 238726 34604
rect 289814 34592 289820 34604
rect 238720 34564 289820 34592
rect 238720 34552 238726 34564
rect 289814 34552 289820 34564
rect 289872 34552 289878 34604
rect 293862 34552 293868 34604
rect 293920 34592 293926 34604
rect 345014 34592 345020 34604
rect 293920 34564 345020 34592
rect 293920 34552 293926 34564
rect 345014 34552 345020 34564
rect 345072 34552 345078 34604
rect 378042 34552 378048 34604
rect 378100 34592 378106 34604
rect 429194 34592 429200 34604
rect 378100 34564 429200 34592
rect 378100 34552 378106 34564
rect 429194 34552 429200 34564
rect 429252 34552 429258 34604
rect 462222 34552 462228 34604
rect 462280 34592 462286 34604
rect 513374 34592 513380 34604
rect 462280 34564 513380 34592
rect 462280 34552 462286 34564
rect 513374 34552 513380 34564
rect 513432 34552 513438 34604
rect 518802 34552 518808 34604
rect 518860 34592 518866 34604
rect 569954 34592 569960 34604
rect 518860 34564 569960 34592
rect 518860 34552 518866 34564
rect 569954 34552 569960 34564
rect 570012 34552 570018 34604
rect 70302 34484 70308 34536
rect 70360 34524 70366 34536
rect 121454 34524 121460 34536
rect 70360 34496 121460 34524
rect 70360 34484 70366 34496
rect 121454 34484 121460 34496
rect 121512 34484 121518 34536
rect 154482 34484 154488 34536
rect 154540 34524 154546 34536
rect 205634 34524 205640 34536
rect 154540 34496 205640 34524
rect 154540 34484 154546 34496
rect 205634 34484 205640 34496
rect 205692 34484 205698 34536
rect 209682 34484 209688 34536
rect 209740 34524 209746 34536
rect 262214 34524 262220 34536
rect 209740 34496 262220 34524
rect 209740 34484 209746 34496
rect 262214 34484 262220 34496
rect 262272 34484 262278 34536
rect 266262 34484 266268 34536
rect 266320 34524 266326 34536
rect 317414 34524 317420 34536
rect 266320 34496 317420 34524
rect 266320 34484 266326 34496
rect 317414 34484 317420 34496
rect 317472 34484 317478 34536
rect 322842 34484 322848 34536
rect 322900 34524 322906 34536
rect 373994 34524 374000 34536
rect 322900 34496 374000 34524
rect 322900 34484 322906 34496
rect 373994 34484 374000 34496
rect 374052 34484 374058 34536
rect 405642 34484 405648 34536
rect 405700 34524 405706 34536
rect 458174 34524 458180 34536
rect 405700 34496 458180 34524
rect 405700 34484 405706 34496
rect 458174 34484 458180 34496
rect 458232 34484 458238 34536
rect 489822 34484 489828 34536
rect 489880 34524 489886 34536
rect 542354 34524 542360 34536
rect 489880 34496 542360 34524
rect 489880 34484 489886 34496
rect 542354 34484 542360 34496
rect 542412 34484 542418 34536
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 12434 33096 12440 33108
rect 7616 33068 12440 33096
rect 7616 33056 7622 33068
rect 12434 33056 12440 33068
rect 12492 33056 12498 33108
rect 63494 27548 63500 27600
rect 63552 27588 63558 27600
rect 68278 27588 68284 27600
rect 63552 27560 68284 27588
rect 63552 27548 63558 27560
rect 68278 27548 68284 27560
rect 68336 27548 68342 27600
rect 259730 21428 259736 21480
rect 259788 21468 259794 21480
rect 260190 21468 260196 21480
rect 259788 21440 260196 21468
rect 259788 21428 259794 21440
rect 260190 21428 260196 21440
rect 260248 21428 260254 21480
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 12434 19292 12440 19304
rect 8996 19264 12440 19292
rect 8996 19252 9002 19264
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 428642 18572 428648 18624
rect 428700 18612 428706 18624
rect 435726 18612 435732 18624
rect 428700 18584 435732 18612
rect 428700 18572 428706 18584
rect 435726 18572 435732 18584
rect 435784 18572 435790 18624
rect 287698 18232 287704 18284
rect 287756 18272 287762 18284
rect 295702 18272 295708 18284
rect 287756 18244 295708 18272
rect 287756 18232 287762 18244
rect 295702 18232 295708 18244
rect 295760 18232 295766 18284
rect 316770 18096 316776 18148
rect 316828 18136 316834 18148
rect 323670 18136 323676 18148
rect 316828 18108 323676 18136
rect 316828 18096 316834 18108
rect 323670 18096 323676 18108
rect 323728 18096 323734 18148
rect 232682 17960 232688 18012
rect 232740 18000 232746 18012
rect 239766 18000 239772 18012
rect 232740 17972 239772 18000
rect 232740 17960 232746 17972
rect 239766 17960 239772 17972
rect 239824 17960 239830 18012
rect 483658 17960 483664 18012
rect 483716 18000 483722 18012
rect 491662 18000 491668 18012
rect 483716 17972 491668 18000
rect 483716 17960 483722 17972
rect 491662 17960 491668 17972
rect 491720 17960 491726 18012
rect 512730 17960 512736 18012
rect 512788 18000 512794 18012
rect 519630 18000 519636 18012
rect 512788 17972 519636 18000
rect 512788 17960 512794 17972
rect 519630 17960 519636 17972
rect 519688 17960 519694 18012
rect 231670 16532 231676 16584
rect 231728 16572 231734 16584
rect 232590 16572 232596 16584
rect 231728 16544 232596 16572
rect 231728 16532 231734 16544
rect 232590 16532 232596 16544
rect 232648 16532 232654 16584
rect 343542 16532 343548 16584
rect 343600 16572 343606 16584
rect 345658 16572 345664 16584
rect 343600 16544 345664 16572
rect 343600 16532 343606 16544
rect 345658 16532 345664 16544
rect 345716 16532 345722 16584
rect 539502 16532 539508 16584
rect 539560 16572 539566 16584
rect 542998 16572 543004 16584
rect 539560 16544 543004 16572
rect 539560 16532 539566 16544
rect 542998 16532 543004 16544
rect 543056 16532 543062 16584
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 16022 13784 16028 13796
rect 6328 13756 16028 13784
rect 6328 13744 6334 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 50154 13744 50160 13796
rect 50212 13784 50218 13796
rect 65518 13784 65524 13796
rect 50212 13756 65524 13784
rect 50212 13744 50218 13756
rect 65518 13744 65524 13756
rect 65576 13744 65582 13796
rect 81986 13744 81992 13796
rect 82044 13784 82050 13796
rect 93118 13784 93124 13796
rect 82044 13756 93124 13784
rect 82044 13744 82050 13756
rect 93118 13744 93124 13756
rect 93176 13744 93182 13796
rect 119338 13744 119344 13796
rect 119396 13784 119402 13796
rect 126238 13784 126244 13796
rect 119396 13756 126244 13784
rect 119396 13744 119402 13756
rect 126238 13744 126244 13756
rect 126296 13744 126302 13796
rect 178678 13744 178684 13796
rect 178736 13784 178742 13796
rect 184014 13784 184020 13796
rect 178736 13756 184020 13784
rect 178736 13744 178742 13756
rect 184014 13744 184020 13756
rect 184072 13744 184078 13796
rect 193674 13744 193680 13796
rect 193732 13784 193738 13796
rect 204898 13784 204904 13796
rect 193732 13756 204904 13784
rect 193732 13744 193738 13756
rect 204898 13744 204904 13756
rect 204956 13744 204962 13796
rect 277670 13744 277676 13796
rect 277728 13784 277734 13796
rect 289078 13784 289084 13796
rect 277728 13756 289084 13784
rect 277728 13744 277734 13756
rect 289078 13744 289084 13756
rect 289136 13744 289142 13796
rect 315666 13744 315672 13796
rect 315724 13784 315730 13796
rect 322198 13784 322204 13796
rect 315724 13756 322204 13784
rect 315724 13744 315730 13756
rect 322198 13744 322204 13756
rect 322256 13744 322262 13796
rect 361666 13744 361672 13796
rect 361724 13784 361730 13796
rect 373258 13784 373264 13796
rect 361724 13756 373264 13784
rect 361724 13744 361730 13756
rect 373258 13744 373264 13756
rect 373316 13744 373322 13796
rect 374638 13744 374644 13796
rect 374696 13784 374702 13796
rect 379698 13784 379704 13796
rect 374696 13756 379704 13784
rect 374696 13744 374702 13756
rect 379698 13744 379704 13756
rect 379756 13744 379762 13796
rect 390002 13744 390008 13796
rect 390060 13784 390066 13796
rect 400858 13784 400864 13796
rect 390060 13756 400864 13784
rect 390060 13744 390066 13756
rect 400858 13744 400864 13756
rect 400916 13744 400922 13796
rect 473998 13744 474004 13796
rect 474056 13784 474062 13796
rect 485038 13784 485044 13796
rect 474056 13756 485044 13784
rect 474056 13744 474062 13756
rect 485038 13744 485044 13756
rect 485096 13744 485102 13796
rect 511350 13744 511356 13796
rect 511408 13784 511414 13796
rect 518158 13784 518164 13796
rect 511408 13756 518164 13784
rect 511408 13744 511414 13756
rect 518158 13744 518164 13756
rect 518216 13744 518222 13796
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 18598 13716 18604 13728
rect 10376 13688 18604 13716
rect 10376 13676 10382 13688
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 53374 13676 53380 13728
rect 53432 13716 53438 13728
rect 60734 13716 60740 13728
rect 53432 13688 60740 13716
rect 53432 13676 53438 13688
rect 60734 13676 60740 13688
rect 60792 13676 60798 13728
rect 109678 13676 109684 13728
rect 109736 13716 109742 13728
rect 120718 13716 120724 13728
rect 109736 13688 120724 13716
rect 109736 13676 109742 13688
rect 120718 13676 120724 13688
rect 120776 13676 120782 13728
rect 137646 13676 137652 13728
rect 137704 13716 137710 13728
rect 148410 13716 148416 13728
rect 137704 13688 148416 13716
rect 137704 13676 137710 13688
rect 148410 13676 148416 13688
rect 148468 13676 148474 13728
rect 306006 13676 306012 13728
rect 306064 13716 306070 13728
rect 316678 13716 316684 13728
rect 306064 13688 316684 13716
rect 306064 13676 306070 13688
rect 316678 13676 316684 13688
rect 316736 13676 316742 13728
rect 333698 13676 333704 13728
rect 333756 13716 333762 13728
rect 344278 13716 344284 13728
rect 333756 13688 344284 13716
rect 333756 13676 333762 13688
rect 344278 13676 344284 13688
rect 344336 13676 344342 13728
rect 417694 13676 417700 13728
rect 417752 13716 417758 13728
rect 428550 13716 428556 13728
rect 417752 13688 428556 13716
rect 417752 13676 417758 13688
rect 428550 13676 428556 13688
rect 428608 13676 428614 13728
rect 445662 13676 445668 13728
rect 445720 13716 445726 13728
rect 456150 13716 456156 13728
rect 445720 13688 456156 13716
rect 445720 13676 445726 13688
rect 456150 13676 456156 13688
rect 456208 13676 456214 13728
rect 3878 13608 3884 13660
rect 3936 13648 3942 13660
rect 59814 13648 59820 13660
rect 3936 13620 59820 13648
rect 3936 13608 3942 13620
rect 59814 13608 59820 13620
rect 59872 13608 59878 13660
rect 64322 13608 64328 13660
rect 64380 13648 64386 13660
rect 557534 13648 557540 13660
rect 64380 13620 557540 13648
rect 64380 13608 64386 13620
rect 557534 13608 557540 13620
rect 557592 13608 557598 13660
rect 7650 13540 7656 13592
rect 7708 13580 7714 13592
rect 25038 13580 25044 13592
rect 7708 13552 25044 13580
rect 7708 13540 7714 13552
rect 25038 13540 25044 13552
rect 25096 13540 25102 13592
rect 46934 13540 46940 13592
rect 46992 13580 46998 13592
rect 490558 13580 490564 13592
rect 46992 13552 490564 13580
rect 46992 13540 46998 13552
rect 490558 13540 490564 13552
rect 490616 13540 490622 13592
rect 501690 13540 501696 13592
rect 501748 13580 501754 13592
rect 512638 13580 512644 13592
rect 501748 13552 512644 13580
rect 501748 13540 501754 13552
rect 512638 13540 512644 13552
rect 512696 13540 512702 13592
rect 518986 13540 518992 13592
rect 519044 13580 519050 13592
rect 547874 13580 547880 13592
rect 519044 13552 547880 13580
rect 519044 13540 519050 13552
rect 547874 13540 547880 13552
rect 547932 13540 547938 13592
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 56594 13512 56600 13524
rect 14516 13484 56600 13512
rect 14516 13472 14522 13484
rect 56594 13472 56600 13484
rect 56652 13472 56658 13524
rect 62758 13472 62764 13524
rect 62816 13512 62822 13524
rect 62816 13484 64874 13512
rect 62816 13472 62822 13484
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 21818 13444 21824 13456
rect 4856 13416 21824 13444
rect 4856 13404 4862 13416
rect 21818 13404 21824 13416
rect 21876 13404 21882 13456
rect 34698 13404 34704 13456
rect 34756 13444 34762 13456
rect 64138 13444 64144 13456
rect 34756 13416 64144 13444
rect 34756 13404 34762 13416
rect 64138 13404 64144 13416
rect 64196 13404 64202 13456
rect 64846 13444 64874 13484
rect 71866 13472 71872 13524
rect 71924 13512 71930 13524
rect 100018 13512 100024 13524
rect 71924 13484 100024 13512
rect 71924 13472 71930 13484
rect 100018 13472 100024 13484
rect 100076 13472 100082 13524
rect 127986 13512 127992 13524
rect 103486 13484 127992 13512
rect 72050 13444 72056 13456
rect 64846 13416 72056 13444
rect 72050 13404 72056 13416
rect 72108 13404 72114 13456
rect 99466 13404 99472 13456
rect 99524 13444 99530 13456
rect 103486 13444 103514 13484
rect 127986 13472 127992 13484
rect 128044 13472 128050 13524
rect 156046 13512 156052 13524
rect 132466 13484 156052 13512
rect 99524 13416 103514 13444
rect 99524 13404 99530 13416
rect 127066 13404 127072 13456
rect 127124 13444 127130 13456
rect 132466 13444 132494 13484
rect 156046 13472 156052 13484
rect 156104 13472 156110 13524
rect 165982 13472 165988 13524
rect 166040 13512 166046 13524
rect 177298 13512 177304 13524
rect 166040 13484 177304 13512
rect 166040 13472 166046 13484
rect 177298 13472 177304 13484
rect 177356 13472 177362 13524
rect 183646 13472 183652 13524
rect 183704 13512 183710 13524
rect 211706 13512 211712 13524
rect 183704 13484 211712 13512
rect 183704 13472 183710 13484
rect 211706 13472 211712 13484
rect 211764 13472 211770 13524
rect 222010 13472 222016 13524
rect 222068 13512 222074 13524
rect 232498 13512 232504 13524
rect 222068 13484 232504 13512
rect 222068 13472 222074 13484
rect 232498 13472 232504 13484
rect 232556 13472 232562 13524
rect 249702 13472 249708 13524
rect 249760 13512 249766 13524
rect 260098 13512 260104 13524
rect 249760 13484 260104 13512
rect 249760 13472 249766 13484
rect 260098 13472 260104 13484
rect 260156 13472 260162 13524
rect 261478 13472 261484 13524
rect 261536 13512 261542 13524
rect 567194 13512 567200 13524
rect 261536 13484 567200 13512
rect 261536 13472 261542 13484
rect 567194 13472 567200 13484
rect 567252 13472 567258 13524
rect 127124 13416 132494 13444
rect 127124 13404 127130 13416
rect 238846 13404 238852 13456
rect 238904 13444 238910 13456
rect 268010 13444 268016 13456
rect 238904 13416 268016 13444
rect 238904 13404 238910 13416
rect 268010 13404 268016 13416
rect 268068 13404 268074 13456
rect 323026 13404 323032 13456
rect 323084 13444 323090 13456
rect 352006 13444 352012 13456
rect 323084 13416 352012 13444
rect 323084 13404 323090 13416
rect 352006 13404 352012 13416
rect 352064 13404 352070 13456
rect 379606 13404 379612 13456
rect 379664 13444 379670 13456
rect 408034 13444 408040 13456
rect 379664 13416 408040 13444
rect 379664 13404 379670 13416
rect 408034 13404 408040 13416
rect 408092 13404 408098 13456
rect 434806 13404 434812 13456
rect 434864 13444 434870 13456
rect 463694 13444 463700 13456
rect 434864 13416 463700 13444
rect 434864 13404 434870 13416
rect 463694 13404 463700 13416
rect 463752 13404 463758 13456
rect 529658 13404 529664 13456
rect 529716 13444 529722 13456
rect 547138 13444 547144 13456
rect 529716 13416 547144 13444
rect 529716 13404 529722 13416
rect 547138 13404 547144 13416
rect 547196 13404 547202 13456
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 31478 13376 31484 13388
rect 4120 13348 31484 13376
rect 4120 13336 4126 13348
rect 31478 13336 31484 13348
rect 31536 13336 31542 13388
rect 40494 13336 40500 13388
rect 40552 13376 40558 13388
rect 567930 13376 567936 13388
rect 40552 13348 567936 13376
rect 40552 13336 40558 13348
rect 567930 13336 567936 13348
rect 567988 13336 567994 13388
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 28258 13308 28264 13320
rect 3844 13280 28264 13308
rect 3844 13268 3850 13280
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 37918 13268 37924 13320
rect 37976 13308 37982 13320
rect 541618 13308 541624 13320
rect 37976 13280 541624 13308
rect 37976 13268 37982 13280
rect 541618 13268 541624 13280
rect 541676 13268 541682 13320
rect 3418 13064 3424 13116
rect 3476 13104 3482 13116
rect 43714 13104 43720 13116
rect 3476 13076 43720 13104
rect 3476 13064 3482 13076
rect 43714 13064 43720 13076
rect 43772 13064 43778 13116
<< via1 >>
rect 68284 700612 68336 700664
rect 105452 700612 105504 700664
rect 64144 700544 64196 700596
rect 170312 700544 170364 700596
rect 36636 700476 36688 700528
rect 300124 700476 300176 700528
rect 64236 700408 64288 700460
rect 364984 700408 365036 700460
rect 65524 700340 65576 700392
rect 429844 700340 429896 700392
rect 36544 700272 36596 700324
rect 559656 700272 559708 700324
rect 490564 699660 490616 699712
rect 494796 699660 494848 699712
rect 25688 686060 25740 686112
rect 71044 686060 71096 686112
rect 212356 686060 212408 686112
rect 232688 686060 232740 686112
rect 296352 686060 296404 686112
rect 316776 686060 316828 686112
rect 408040 686060 408092 686112
rect 428648 686060 428700 686112
rect 492036 686060 492088 686112
rect 512736 686060 512788 686112
rect 36912 685992 36964 686044
rect 53656 685992 53708 686044
rect 64328 685992 64380 686044
rect 81440 685992 81492 686044
rect 148416 685992 148468 686044
rect 165712 685992 165764 686044
rect 175464 685992 175516 686044
rect 193680 685992 193732 686044
rect 203524 685992 203576 686044
rect 221372 685992 221424 686044
rect 260196 685992 260248 686044
rect 277676 685992 277728 686044
rect 287520 685992 287572 686044
rect 305368 685992 305420 686044
rect 345664 685992 345716 686044
rect 361672 685992 361724 686044
rect 371516 685992 371568 686044
rect 389364 685992 389416 686044
rect 399484 685992 399536 686044
rect 417700 685992 417752 686044
rect 456156 685992 456208 686044
rect 473360 685992 473412 686044
rect 483480 685992 483532 686044
rect 501696 685992 501748 686044
rect 36820 685924 36872 685976
rect 63316 685924 63368 685976
rect 66904 685924 66956 685976
rect 91100 685924 91152 685976
rect 91468 685924 91520 685976
rect 109684 685924 109736 685976
rect 119436 685924 119488 685976
rect 137652 685924 137704 685976
rect 156328 685924 156380 685976
rect 178684 685924 178736 685976
rect 232504 685924 232556 685976
rect 249708 685924 249760 685976
rect 268016 685924 268068 685976
rect 287704 685924 287756 685976
rect 315488 685924 315540 685976
rect 333704 685924 333756 685976
rect 352012 685924 352064 685976
rect 374644 685924 374696 685976
rect 428464 685924 428516 685976
rect 445668 685924 445720 685976
rect 464344 685924 464396 685976
rect 483664 685924 483716 685976
rect 511448 685924 511500 685976
rect 529664 685924 529716 685976
rect 543004 685924 543056 685976
rect 557540 685924 557592 685976
rect 94504 685856 94556 685908
rect 119344 685856 119396 685908
rect 120724 685856 120776 685908
rect 147312 685856 147364 685908
rect 148324 685856 148376 685908
rect 175372 685856 175424 685908
rect 177304 685856 177356 685908
rect 203340 685856 203392 685908
rect 204904 685856 204956 685908
rect 231032 685856 231084 685908
rect 232596 685856 232648 685908
rect 259368 685856 259420 685908
rect 260104 685856 260156 685908
rect 287336 685856 287388 685908
rect 289084 685856 289136 685908
rect 315028 685856 315080 685908
rect 316684 685856 316736 685908
rect 343364 685856 343416 685908
rect 344284 685856 344336 685908
rect 371332 685856 371384 685908
rect 373264 685856 373316 685908
rect 399024 685856 399076 685908
rect 400864 685856 400916 685908
rect 427360 685856 427412 685908
rect 428556 685856 428608 685908
rect 455328 685856 455380 685908
rect 456064 685856 456116 685908
rect 483020 685856 483072 685908
rect 485044 685856 485096 685908
rect 511356 685856 511408 685908
rect 512644 685856 512696 685908
rect 539324 685856 539376 685908
rect 540244 685856 540296 685908
rect 567200 685856 567252 685908
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 182088 683204 182140 683256
rect 233240 683204 233292 683256
rect 378048 683204 378100 683256
rect 429200 683204 429252 683256
rect 35624 683136 35676 683188
rect 36728 683136 36780 683188
rect 42708 683136 42760 683188
rect 93860 683136 93912 683188
rect 97908 683136 97960 683188
rect 149060 683136 149112 683188
rect 154488 683136 154540 683188
rect 205640 683136 205692 683188
rect 238668 683136 238720 683188
rect 289820 683136 289872 683188
rect 293868 683136 293920 683188
rect 345020 683136 345072 683188
rect 350448 683136 350500 683188
rect 401600 683136 401652 683188
rect 434628 683136 434680 683188
rect 485780 683136 485832 683188
rect 489828 683136 489880 683188
rect 542360 683136 542412 683188
rect 541624 673820 541676 673872
rect 545120 673820 545172 673872
rect 567844 670692 567896 670744
rect 580172 670692 580224 670744
rect 63592 668720 63644 668772
rect 64328 668720 64380 668772
rect 147680 668720 147732 668772
rect 148416 668720 148468 668772
rect 259736 668720 259788 668772
rect 260196 668720 260248 668772
rect 455696 668720 455748 668772
rect 456156 668720 456208 668772
rect 428648 665796 428700 665848
rect 435732 665796 435784 665848
rect 287704 665456 287756 665508
rect 295708 665456 295760 665508
rect 316776 665456 316828 665508
rect 323676 665456 323728 665508
rect 232688 665252 232740 665304
rect 239772 665252 239824 665304
rect 483664 665252 483716 665304
rect 491668 665252 491720 665304
rect 512736 665252 512788 665304
rect 519636 665252 519688 665304
rect 13728 665116 13780 665168
rect 66260 665116 66312 665168
rect 70308 665116 70360 665168
rect 121460 665116 121512 665168
rect 126888 665116 126940 665168
rect 178040 665116 178092 665168
rect 209688 665116 209740 665168
rect 262220 665116 262272 665168
rect 266268 665116 266320 665168
rect 317420 665116 317472 665168
rect 322848 665116 322900 665168
rect 374000 665116 374052 665168
rect 405648 665116 405700 665168
rect 458180 665116 458232 665168
rect 462228 665116 462280 665168
rect 513380 665116 513432 665168
rect 518808 665116 518860 665168
rect 569960 665116 570012 665168
rect 35624 665048 35676 665100
rect 36912 665048 36964 665100
rect 343548 665048 343600 665100
rect 345664 665048 345716 665100
rect 71872 662328 71924 662380
rect 100024 662328 100076 662380
rect 25688 662260 25740 662312
rect 36820 662260 36872 662312
rect 42892 662260 42944 662312
rect 15200 662192 15252 662244
rect 43628 662192 43680 662244
rect 53748 662260 53800 662312
rect 66904 662260 66956 662312
rect 81992 662260 82044 662312
rect 94504 662260 94556 662312
rect 99472 662260 99524 662312
rect 127716 662328 127768 662380
rect 165988 662328 166040 662380
rect 177304 662328 177356 662380
rect 178684 662328 178736 662380
rect 184020 662328 184072 662380
rect 109684 662260 109736 662312
rect 120724 662260 120776 662312
rect 137928 662260 137980 662312
rect 148324 662260 148376 662312
rect 183652 662260 183704 662312
rect 211712 662328 211764 662380
rect 277676 662328 277728 662380
rect 289084 662328 289136 662380
rect 306012 662328 306064 662380
rect 316684 662328 316736 662380
rect 361672 662328 361724 662380
rect 373264 662328 373316 662380
rect 374644 662328 374696 662380
rect 379704 662328 379756 662380
rect 193680 662260 193732 662312
rect 204904 662260 204956 662312
rect 222016 662260 222068 662312
rect 232596 662260 232648 662312
rect 249616 662260 249668 662312
rect 260104 662260 260156 662312
rect 333888 662260 333940 662312
rect 344284 662260 344336 662312
rect 379612 662260 379664 662312
rect 408040 662328 408092 662380
rect 474004 662328 474056 662380
rect 485044 662328 485096 662380
rect 501696 662328 501748 662380
rect 512644 662328 512696 662380
rect 518992 662328 519044 662380
rect 547880 662328 547932 662380
rect 390008 662260 390060 662312
rect 400864 662260 400916 662312
rect 417700 662260 417752 662312
rect 428556 662260 428608 662312
rect 445668 662260 445720 662312
rect 456064 662260 456116 662312
rect 539324 662260 539376 662312
rect 543004 662260 543056 662312
rect 71964 662192 72016 662244
rect 127072 662192 127124 662244
rect 155960 662192 156012 662244
rect 238852 662192 238904 662244
rect 268016 662192 268068 662244
rect 323032 662192 323084 662244
rect 352012 662192 352064 662244
rect 434812 662192 434864 662244
rect 463792 662192 463844 662244
rect 529664 662192 529716 662244
rect 540244 662192 540296 662244
rect 16028 658928 16080 658980
rect 547880 658928 547932 658980
rect 25688 658452 25740 658504
rect 66904 658452 66956 658504
rect 212356 658452 212408 658504
rect 232688 658452 232740 658504
rect 296352 658452 296404 658504
rect 316776 658452 316828 658504
rect 408040 658452 408092 658504
rect 428648 658452 428700 658504
rect 492036 658452 492088 658504
rect 512736 658452 512788 658504
rect 37004 658384 37056 658436
rect 53656 658384 53708 658436
rect 148324 658384 148376 658436
rect 165712 658384 165764 658436
rect 175464 658384 175516 658436
rect 193680 658384 193732 658436
rect 203524 658384 203576 658436
rect 221372 658384 221424 658436
rect 260196 658384 260248 658436
rect 277676 658384 277728 658436
rect 287520 658384 287572 658436
rect 305368 658384 305420 658436
rect 345664 658384 345716 658436
rect 361672 658384 361724 658436
rect 371516 658384 371568 658436
rect 389364 658384 389416 658436
rect 399484 658384 399536 658436
rect 417700 658384 417752 658436
rect 456064 658384 456116 658436
rect 473360 658384 473412 658436
rect 483480 658384 483532 658436
rect 501696 658384 501748 658436
rect 36912 658316 36964 658368
rect 63316 658316 63368 658368
rect 64328 658316 64380 658368
rect 81440 658316 81492 658368
rect 91468 658316 91520 658368
rect 109684 658316 109736 658368
rect 119436 658316 119488 658368
rect 137652 658316 137704 658368
rect 156328 658316 156380 658368
rect 178684 658316 178736 658368
rect 232596 658316 232648 658368
rect 249708 658316 249760 658368
rect 268016 658316 268068 658368
rect 287704 658316 287756 658368
rect 315488 658316 315540 658368
rect 333704 658316 333756 658368
rect 352012 658316 352064 658368
rect 374644 658316 374696 658368
rect 428464 658316 428516 658368
rect 445668 658316 445720 658368
rect 464344 658316 464396 658368
rect 483664 658316 483716 658368
rect 511448 658316 511500 658368
rect 529664 658316 529716 658368
rect 543004 658316 543056 658368
rect 557540 658316 557592 658368
rect 69664 658248 69716 658300
rect 91100 658248 91152 658300
rect 94504 658248 94556 658300
rect 119344 658248 119396 658300
rect 120724 658248 120776 658300
rect 147312 658248 147364 658300
rect 148416 658248 148468 658300
rect 175372 658248 175424 658300
rect 177304 658248 177356 658300
rect 203340 658248 203392 658300
rect 204904 658248 204956 658300
rect 231032 658248 231084 658300
rect 232504 658248 232556 658300
rect 259368 658248 259420 658300
rect 260104 658248 260156 658300
rect 287336 658248 287388 658300
rect 289084 658248 289136 658300
rect 315028 658248 315080 658300
rect 316684 658248 316736 658300
rect 343364 658248 343416 658300
rect 344284 658248 344336 658300
rect 371332 658248 371384 658300
rect 373264 658248 373316 658300
rect 399024 658248 399076 658300
rect 400864 658248 400916 658300
rect 427360 658248 427412 658300
rect 428556 658248 428608 658300
rect 455328 658248 455380 658300
rect 456156 658248 456208 658300
rect 483020 658248 483072 658300
rect 485044 658248 485096 658300
rect 511356 658248 511408 658300
rect 512644 658248 512696 658300
rect 539324 658248 539376 658300
rect 540244 658248 540296 658300
rect 567200 658248 567252 658300
rect 37924 657500 37976 657552
rect 545764 657500 545816 657552
rect 35624 656888 35676 656940
rect 36820 656888 36872 656940
rect 183560 655664 183612 655716
rect 233240 655664 233292 655716
rect 378048 655664 378100 655716
rect 429200 655664 429252 655716
rect 463700 655664 463752 655716
rect 513380 655664 513432 655716
rect 42708 655596 42760 655648
rect 93860 655596 93912 655648
rect 97908 655596 97960 655648
rect 149060 655596 149112 655648
rect 154488 655596 154540 655648
rect 205640 655596 205692 655648
rect 238668 655596 238720 655648
rect 289820 655596 289872 655648
rect 293868 655596 293920 655648
rect 345020 655596 345072 655648
rect 350448 655596 350500 655648
rect 401600 655596 401652 655648
rect 434628 655596 434680 655648
rect 485780 655596 485832 655648
rect 518808 655596 518860 655648
rect 569960 655596 570012 655648
rect 13728 655528 13780 655580
rect 66260 655528 66312 655580
rect 70308 655528 70360 655580
rect 121460 655528 121512 655580
rect 126888 655528 126940 655580
rect 178040 655528 178092 655580
rect 209688 655528 209740 655580
rect 262220 655528 262272 655580
rect 266268 655528 266320 655580
rect 317420 655528 317472 655580
rect 322848 655528 322900 655580
rect 374000 655528 374052 655580
rect 405648 655528 405700 655580
rect 458180 655528 458232 655580
rect 489828 655528 489880 655580
rect 542360 655528 542412 655580
rect 182088 654032 182140 654084
rect 183560 654032 183612 654084
rect 462228 654032 462280 654084
rect 463700 654032 463752 654084
rect 63592 640772 63644 640824
rect 64328 640772 64380 640824
rect 259736 640772 259788 640824
rect 260196 640772 260248 640824
rect 287704 639752 287756 639804
rect 295708 639752 295760 639804
rect 428648 639548 428700 639600
rect 435732 639548 435784 639600
rect 232688 639344 232740 639396
rect 239772 639344 239824 639396
rect 316776 639344 316828 639396
rect 323676 639344 323728 639396
rect 483664 639344 483716 639396
rect 491668 639344 491720 639396
rect 512736 639072 512788 639124
rect 519636 639072 519688 639124
rect 35624 637508 35676 637560
rect 37004 637508 37056 637560
rect 343640 637508 343692 637560
rect 345664 637508 345716 637560
rect 25688 634720 25740 634772
rect 36912 634720 36964 634772
rect 178684 634720 178736 634772
rect 184020 634720 184072 634772
rect 231584 634720 231636 634772
rect 232596 634720 232648 634772
rect 374644 634720 374696 634772
rect 379704 634720 379756 634772
rect 539324 634720 539376 634772
rect 543004 634720 543056 634772
rect 15200 634652 15252 634704
rect 43996 634652 44048 634704
rect 71044 634652 71096 634704
rect 567200 634652 567252 634704
rect 53656 634584 53708 634636
rect 69664 634584 69716 634636
rect 71872 634584 71924 634636
rect 100024 634584 100076 634636
rect 42892 634516 42944 634568
rect 71964 634516 72016 634568
rect 81992 634516 82044 634568
rect 94504 634516 94556 634568
rect 99472 634516 99524 634568
rect 127992 634584 128044 634636
rect 109684 634516 109736 634568
rect 120724 634516 120776 634568
rect 127072 634516 127124 634568
rect 155960 634584 156012 634636
rect 165988 634584 166040 634636
rect 177304 634584 177356 634636
rect 183652 634584 183704 634636
rect 211712 634584 211764 634636
rect 221924 634584 221976 634636
rect 232504 634584 232556 634636
rect 238852 634584 238904 634636
rect 268016 634584 268068 634636
rect 277676 634584 277728 634636
rect 289084 634584 289136 634636
rect 306012 634584 306064 634636
rect 316684 634584 316736 634636
rect 323032 634584 323084 634636
rect 352012 634584 352064 634636
rect 361672 634584 361724 634636
rect 373264 634584 373316 634636
rect 379612 634584 379664 634636
rect 408040 634584 408092 634636
rect 417700 634584 417752 634636
rect 428556 634584 428608 634636
rect 434812 634584 434864 634636
rect 463792 634584 463844 634636
rect 474004 634584 474056 634636
rect 485044 634584 485096 634636
rect 501696 634584 501748 634636
rect 512644 634584 512696 634636
rect 518992 634584 519044 634636
rect 547880 634584 547932 634636
rect 137652 634516 137704 634568
rect 148416 634516 148468 634568
rect 193680 634516 193732 634568
rect 204904 634516 204956 634568
rect 249708 634516 249760 634568
rect 260104 634516 260156 634568
rect 333704 634516 333756 634568
rect 344284 634516 344336 634568
rect 390008 634516 390060 634568
rect 400864 634516 400916 634568
rect 445668 634516 445720 634568
rect 456156 634516 456208 634568
rect 529664 634516 529716 634568
rect 540244 634516 540296 634568
rect 36728 634448 36780 634500
rect 557540 634448 557592 634500
rect 16028 632680 16080 632732
rect 547880 632680 547932 632732
rect 25688 632272 25740 632324
rect 71044 632272 71096 632324
rect 212356 632272 212408 632324
rect 232688 632272 232740 632324
rect 408040 632272 408092 632324
rect 428648 632272 428700 632324
rect 492036 632272 492088 632324
rect 512736 632272 512788 632324
rect 37004 632204 37056 632256
rect 53656 632204 53708 632256
rect 148324 632204 148376 632256
rect 165712 632204 165764 632256
rect 175464 632204 175516 632256
rect 193680 632204 193732 632256
rect 203524 632204 203576 632256
rect 221372 632204 221424 632256
rect 260104 632204 260156 632256
rect 277676 632204 277728 632256
rect 287520 632204 287572 632256
rect 305368 632204 305420 632256
rect 315488 632204 315540 632256
rect 333704 632204 333756 632256
rect 345664 632204 345716 632256
rect 361672 632204 361724 632256
rect 371516 632204 371568 632256
rect 389364 632204 389416 632256
rect 399484 632204 399536 632256
rect 417700 632204 417752 632256
rect 456156 632204 456208 632256
rect 473360 632204 473412 632256
rect 483480 632204 483532 632256
rect 501696 632204 501748 632256
rect 36912 632136 36964 632188
rect 63316 632136 63368 632188
rect 64328 632136 64380 632188
rect 81440 632136 81492 632188
rect 91468 632136 91520 632188
rect 109684 632136 109736 632188
rect 119436 632136 119488 632188
rect 137652 632136 137704 632188
rect 156328 632136 156380 632188
rect 178684 632136 178736 632188
rect 232596 632136 232648 632188
rect 249708 632136 249760 632188
rect 268016 632136 268068 632188
rect 287704 632136 287756 632188
rect 296352 632136 296404 632188
rect 316776 632136 316828 632188
rect 352012 632136 352064 632188
rect 374644 632136 374696 632188
rect 428464 632136 428516 632188
rect 445668 632136 445720 632188
rect 464344 632136 464396 632188
rect 483664 632136 483716 632188
rect 511448 632136 511500 632188
rect 529664 632136 529716 632188
rect 543004 632136 543056 632188
rect 557540 632136 557592 632188
rect 3148 632068 3200 632120
rect 6184 632068 6236 632120
rect 69664 632068 69716 632120
rect 91100 632068 91152 632120
rect 95884 632068 95936 632120
rect 119344 632068 119396 632120
rect 120724 632068 120776 632120
rect 147312 632068 147364 632120
rect 148416 632068 148468 632120
rect 175372 632068 175424 632120
rect 177304 632068 177356 632120
rect 203340 632068 203392 632120
rect 204904 632068 204956 632120
rect 231032 632068 231084 632120
rect 232504 632068 232556 632120
rect 259368 632068 259420 632120
rect 260196 632068 260248 632120
rect 287336 632068 287388 632120
rect 289084 632068 289136 632120
rect 315028 632068 315080 632120
rect 316684 632068 316736 632120
rect 343364 632068 343416 632120
rect 344284 632068 344336 632120
rect 371332 632068 371384 632120
rect 373264 632068 373316 632120
rect 399024 632068 399076 632120
rect 400864 632068 400916 632120
rect 427360 632068 427412 632120
rect 428556 632068 428608 632120
rect 455328 632068 455380 632120
rect 456064 632068 456116 632120
rect 483020 632068 483072 632120
rect 485044 632068 485096 632120
rect 511356 632068 511408 632120
rect 512644 632068 512696 632120
rect 539324 632068 539376 632120
rect 540244 632068 540296 632120
rect 567200 632068 567252 632120
rect 37924 629892 37976 629944
rect 545764 629892 545816 629944
rect 35624 629280 35676 629332
rect 36728 629280 36780 629332
rect 567936 616836 567988 616888
rect 580172 616836 580224 616888
rect 63592 612756 63644 612808
rect 64328 612756 64380 612808
rect 455696 612756 455748 612808
rect 456156 612756 456208 612808
rect 316776 612008 316828 612060
rect 323676 612008 323728 612060
rect 428648 612008 428700 612060
rect 435732 612008 435784 612060
rect 232688 611940 232740 611992
rect 239772 611940 239824 611992
rect 287704 611872 287756 611924
rect 295708 611872 295760 611924
rect 483664 611736 483716 611788
rect 491668 611736 491720 611788
rect 512736 611736 512788 611788
rect 519636 611736 519688 611788
rect 13728 611260 13780 611312
rect 66260 611260 66312 611312
rect 70308 611260 70360 611312
rect 121460 611260 121512 611312
rect 126888 611260 126940 611312
rect 178040 611260 178092 611312
rect 209688 611260 209740 611312
rect 262220 611260 262272 611312
rect 266268 611260 266320 611312
rect 317420 611260 317472 611312
rect 322848 611260 322900 611312
rect 374000 611260 374052 611312
rect 405648 611260 405700 611312
rect 458180 611260 458232 611312
rect 489828 611260 489880 611312
rect 542360 611260 542412 611312
rect 35624 611192 35676 611244
rect 37004 611192 37056 611244
rect 42708 611192 42760 611244
rect 93860 611192 93912 611244
rect 97908 611192 97960 611244
rect 149060 611192 149112 611244
rect 154488 611192 154540 611244
rect 205640 611192 205692 611244
rect 231676 611192 231728 611244
rect 232596 611192 232648 611244
rect 238668 611192 238720 611244
rect 289820 611192 289872 611244
rect 293868 611192 293920 611244
rect 345020 611192 345072 611244
rect 350448 611192 350500 611244
rect 401600 611192 401652 611244
rect 462228 611192 462280 611244
rect 513380 611192 513432 611244
rect 518808 611192 518860 611244
rect 569960 611192 570012 611244
rect 182088 611124 182140 611176
rect 233240 611124 233292 611176
rect 378048 611124 378100 611176
rect 429200 611124 429252 611176
rect 434628 611124 434680 611176
rect 485780 611124 485832 611176
rect 15200 608472 15252 608524
rect 43996 608472 44048 608524
rect 25688 608404 25740 608456
rect 36912 608404 36964 608456
rect 42892 608404 42944 608456
rect 72056 608540 72108 608592
rect 178684 608540 178736 608592
rect 184020 608540 184072 608592
rect 343364 608540 343416 608592
rect 345664 608540 345716 608592
rect 374644 608540 374696 608592
rect 379704 608540 379756 608592
rect 539324 608540 539376 608592
rect 543004 608540 543056 608592
rect 66904 608472 66956 608524
rect 567200 608472 567252 608524
rect 71872 608404 71924 608456
rect 100024 608404 100076 608456
rect 53656 608336 53708 608388
rect 69664 608336 69716 608388
rect 81992 608336 82044 608388
rect 95884 608336 95936 608388
rect 99472 608336 99524 608388
rect 127992 608404 128044 608456
rect 109684 608336 109736 608388
rect 120724 608336 120776 608388
rect 127072 608336 127124 608388
rect 156052 608404 156104 608456
rect 165988 608404 166040 608456
rect 177304 608404 177356 608456
rect 183652 608404 183704 608456
rect 211712 608404 211764 608456
rect 222016 608404 222068 608456
rect 232504 608404 232556 608456
rect 238852 608404 238904 608456
rect 268016 608404 268068 608456
rect 277676 608404 277728 608456
rect 289084 608404 289136 608456
rect 306012 608404 306064 608456
rect 316684 608404 316736 608456
rect 323032 608404 323084 608456
rect 352012 608404 352064 608456
rect 361672 608404 361724 608456
rect 373264 608404 373316 608456
rect 379612 608404 379664 608456
rect 408040 608404 408092 608456
rect 417700 608404 417752 608456
rect 428556 608404 428608 608456
rect 434812 608404 434864 608456
rect 463700 608404 463752 608456
rect 474004 608404 474056 608456
rect 485044 608404 485096 608456
rect 501696 608404 501748 608456
rect 512644 608404 512696 608456
rect 518992 608404 519044 608456
rect 547880 608404 547932 608456
rect 137652 608336 137704 608388
rect 148416 608336 148468 608388
rect 193680 608336 193732 608388
rect 204904 608336 204956 608388
rect 249708 608336 249760 608388
rect 260196 608336 260248 608388
rect 333704 608336 333756 608388
rect 344284 608336 344336 608388
rect 390008 608336 390060 608388
rect 400864 608336 400916 608388
rect 445668 608336 445720 608388
rect 456064 608336 456116 608388
rect 529664 608336 529716 608388
rect 540244 608336 540296 608388
rect 36820 608268 36872 608320
rect 557540 608268 557592 608320
rect 15292 605072 15344 605124
rect 547880 605072 547932 605124
rect 25688 604732 25740 604784
rect 261484 604732 261536 604784
rect 119436 604664 119488 604716
rect 137652 604664 137704 604716
rect 148324 604664 148376 604716
rect 165712 604664 165764 604716
rect 175464 604664 175516 604716
rect 193680 604664 193732 604716
rect 203524 604664 203576 604716
rect 221372 604664 221424 604716
rect 408040 604664 408092 604716
rect 428648 604664 428700 604716
rect 492036 604664 492088 604716
rect 512736 604664 512788 604716
rect 37004 604596 37056 604648
rect 53656 604596 53708 604648
rect 64328 604596 64380 604648
rect 81440 604596 81492 604648
rect 91468 604596 91520 604648
rect 109684 604596 109736 604648
rect 127992 604596 128044 604648
rect 148508 604596 148560 604648
rect 156328 604596 156380 604648
rect 178684 604596 178736 604648
rect 232504 604596 232556 604648
rect 249708 604596 249760 604648
rect 260196 604596 260248 604648
rect 277676 604596 277728 604648
rect 287520 604596 287572 604648
rect 305368 604596 305420 604648
rect 315488 604596 315540 604648
rect 333704 604596 333756 604648
rect 345664 604596 345716 604648
rect 361672 604596 361724 604648
rect 371516 604596 371568 604648
rect 389364 604596 389416 604648
rect 399484 604596 399536 604648
rect 417700 604596 417752 604648
rect 456064 604596 456116 604648
rect 473360 604596 473412 604648
rect 483480 604596 483532 604648
rect 501696 604596 501748 604648
rect 36912 604528 36964 604580
rect 63316 604528 63368 604580
rect 66904 604528 66956 604580
rect 91100 604528 91152 604580
rect 94504 604528 94556 604580
rect 119344 604528 119396 604580
rect 120724 604528 120776 604580
rect 147312 604528 147364 604580
rect 148416 604528 148468 604580
rect 175372 604528 175424 604580
rect 177304 604528 177356 604580
rect 203340 604528 203392 604580
rect 204904 604528 204956 604580
rect 231032 604528 231084 604580
rect 232596 604528 232648 604580
rect 259368 604528 259420 604580
rect 268016 604528 268068 604580
rect 287704 604528 287756 604580
rect 296352 604528 296404 604580
rect 316776 604528 316828 604580
rect 352012 604528 352064 604580
rect 374644 604528 374696 604580
rect 428556 604528 428608 604580
rect 445668 604528 445720 604580
rect 464344 604528 464396 604580
rect 483664 604528 483716 604580
rect 511448 604528 511500 604580
rect 529664 604528 529716 604580
rect 543004 604528 543056 604580
rect 557540 604528 557592 604580
rect 212356 604460 212408 604512
rect 232688 604460 232740 604512
rect 260104 604460 260156 604512
rect 287336 604460 287388 604512
rect 289084 604460 289136 604512
rect 315028 604460 315080 604512
rect 316684 604460 316736 604512
rect 343364 604460 343416 604512
rect 344284 604460 344336 604512
rect 371332 604460 371384 604512
rect 373264 604460 373316 604512
rect 399024 604460 399076 604512
rect 400864 604460 400916 604512
rect 427360 604460 427412 604512
rect 428464 604460 428516 604512
rect 455328 604460 455380 604512
rect 456156 604460 456208 604512
rect 483020 604460 483072 604512
rect 485044 604460 485096 604512
rect 511356 604460 511408 604512
rect 512644 604460 512696 604512
rect 539324 604460 539376 604512
rect 540244 604460 540296 604512
rect 567200 604460 567252 604512
rect 37924 602352 37976 602404
rect 545764 602352 545816 602404
rect 35624 601672 35676 601724
rect 36820 601672 36872 601724
rect 259736 584740 259788 584792
rect 260196 584740 260248 584792
rect 148508 584400 148560 584452
rect 155868 584400 155920 584452
rect 232688 584400 232740 584452
rect 239772 584400 239824 584452
rect 428648 584400 428700 584452
rect 435732 584400 435784 584452
rect 316776 584264 316828 584316
rect 323860 584264 323912 584316
rect 512736 584264 512788 584316
rect 519636 584264 519688 584316
rect 287704 584128 287756 584180
rect 295708 584128 295760 584180
rect 483664 584128 483716 584180
rect 491668 584128 491720 584180
rect 13728 583652 13780 583704
rect 35624 583584 35676 583636
rect 37004 583584 37056 583636
rect 42708 583584 42760 583636
rect 63592 583652 63644 583704
rect 64328 583652 64380 583704
rect 70308 583652 70360 583704
rect 121460 583652 121512 583704
rect 126888 583652 126940 583704
rect 178040 583652 178092 583704
rect 209688 583652 209740 583704
rect 262220 583652 262272 583704
rect 266268 583652 266320 583704
rect 317420 583652 317472 583704
rect 322848 583652 322900 583704
rect 374000 583652 374052 583704
rect 405648 583652 405700 583704
rect 458180 583652 458232 583704
rect 489828 583652 489880 583704
rect 542360 583652 542412 583704
rect 66260 583516 66312 583568
rect 93860 583584 93912 583636
rect 97908 583584 97960 583636
rect 149060 583584 149112 583636
rect 154488 583584 154540 583636
rect 205640 583584 205692 583636
rect 238668 583584 238720 583636
rect 289820 583584 289872 583636
rect 293868 583584 293920 583636
rect 182088 583516 182140 583568
rect 233240 583516 233292 583568
rect 343640 583584 343692 583636
rect 345664 583584 345716 583636
rect 350448 583584 350500 583636
rect 401600 583584 401652 583636
rect 427728 583584 427780 583636
rect 428556 583584 428608 583636
rect 434628 583584 434680 583636
rect 485780 583584 485832 583636
rect 518808 583584 518860 583636
rect 569960 583584 570012 583636
rect 345020 583516 345072 583568
rect 378048 583516 378100 583568
rect 429200 583516 429252 583568
rect 462228 583516 462280 583568
rect 513380 583516 513432 583568
rect 539508 583516 539560 583568
rect 543004 583516 543056 583568
rect 178684 580932 178736 580984
rect 184020 580932 184072 580984
rect 374644 580932 374696 580984
rect 379704 580932 379756 580984
rect 15200 580864 15252 580916
rect 43996 580864 44048 580916
rect 71044 580864 71096 580916
rect 567200 580864 567252 580916
rect 25688 580796 25740 580848
rect 36912 580796 36964 580848
rect 53656 580796 53708 580848
rect 66904 580796 66956 580848
rect 71872 580796 71924 580848
rect 100024 580796 100076 580848
rect 42892 580728 42944 580780
rect 72056 580728 72108 580780
rect 81992 580728 82044 580780
rect 94504 580728 94556 580780
rect 99472 580728 99524 580780
rect 127992 580796 128044 580848
rect 137652 580796 137704 580848
rect 148416 580796 148468 580848
rect 165988 580796 166040 580848
rect 177304 580796 177356 580848
rect 183652 580796 183704 580848
rect 211712 580796 211764 580848
rect 222016 580796 222068 580848
rect 232596 580796 232648 580848
rect 238852 580796 238904 580848
rect 268016 580796 268068 580848
rect 277676 580796 277728 580848
rect 289084 580796 289136 580848
rect 306012 580796 306064 580848
rect 316684 580796 316736 580848
rect 323032 580796 323084 580848
rect 352012 580796 352064 580848
rect 361672 580796 361724 580848
rect 373264 580796 373316 580848
rect 379612 580796 379664 580848
rect 408040 580796 408092 580848
rect 417700 580796 417752 580848
rect 428464 580796 428516 580848
rect 434812 580796 434864 580848
rect 463700 580796 463752 580848
rect 474004 580796 474056 580848
rect 485044 580796 485096 580848
rect 501696 580796 501748 580848
rect 512644 580796 512696 580848
rect 518992 580796 519044 580848
rect 547880 580796 547932 580848
rect 109684 580728 109736 580780
rect 120724 580728 120776 580780
rect 193680 580728 193732 580780
rect 204904 580728 204956 580780
rect 249708 580728 249760 580780
rect 260104 580728 260156 580780
rect 333704 580728 333756 580780
rect 344284 580728 344336 580780
rect 390008 580728 390060 580780
rect 400864 580728 400916 580780
rect 445668 580728 445720 580780
rect 456156 580728 456208 580780
rect 529664 580728 529716 580780
rect 540244 580728 540296 580780
rect 36728 580660 36780 580712
rect 557540 580660 557592 580712
rect 3240 579708 3292 579760
rect 7564 579708 7616 579760
rect 16028 578892 16080 578944
rect 547880 578892 547932 578944
rect 25688 578416 25740 578468
rect 71044 578416 71096 578468
rect 296352 578416 296404 578468
rect 316776 578416 316828 578468
rect 408040 578416 408092 578468
rect 428648 578416 428700 578468
rect 492036 578416 492088 578468
rect 512736 578416 512788 578468
rect 36912 578348 36964 578400
rect 53656 578348 53708 578400
rect 148416 578348 148468 578400
rect 165620 578348 165672 578400
rect 175464 578348 175516 578400
rect 193680 578348 193732 578400
rect 203524 578348 203576 578400
rect 221372 578348 221424 578400
rect 232504 578348 232556 578400
rect 249708 578348 249760 578400
rect 260196 578348 260248 578400
rect 277676 578348 277728 578400
rect 287520 578348 287572 578400
rect 305368 578348 305420 578400
rect 345664 578348 345716 578400
rect 361672 578348 361724 578400
rect 371516 578348 371568 578400
rect 389364 578348 389416 578400
rect 399484 578348 399536 578400
rect 417700 578348 417752 578400
rect 456156 578348 456208 578400
rect 473544 578348 473596 578400
rect 483480 578348 483532 578400
rect 501696 578348 501748 578400
rect 37004 578280 37056 578332
rect 63316 578280 63368 578332
rect 64328 578280 64380 578332
rect 81440 578280 81492 578332
rect 91468 578280 91520 578332
rect 109684 578280 109736 578332
rect 119436 578280 119488 578332
rect 137652 578280 137704 578332
rect 156328 578280 156380 578332
rect 178684 578280 178736 578332
rect 212264 578280 212316 578332
rect 232688 578280 232740 578332
rect 268016 578280 268068 578332
rect 287704 578280 287756 578332
rect 315488 578280 315540 578332
rect 333704 578280 333756 578332
rect 352012 578280 352064 578332
rect 374644 578280 374696 578332
rect 428464 578280 428516 578332
rect 445668 578280 445720 578332
rect 464344 578280 464396 578332
rect 483664 578280 483716 578332
rect 511448 578280 511500 578332
rect 529664 578280 529716 578332
rect 543004 578280 543056 578332
rect 557540 578280 557592 578332
rect 69664 578212 69716 578264
rect 91100 578212 91152 578264
rect 94504 578212 94556 578264
rect 119344 578212 119396 578264
rect 120724 578212 120776 578264
rect 147312 578212 147364 578264
rect 148324 578212 148376 578264
rect 175280 578212 175332 578264
rect 177304 578212 177356 578264
rect 203340 578212 203392 578264
rect 204904 578212 204956 578264
rect 231032 578212 231084 578264
rect 232596 578212 232648 578264
rect 259368 578212 259420 578264
rect 260104 578212 260156 578264
rect 287336 578212 287388 578264
rect 289084 578212 289136 578264
rect 315028 578212 315080 578264
rect 316684 578212 316736 578264
rect 343364 578212 343416 578264
rect 344284 578212 344336 578264
rect 371332 578212 371384 578264
rect 373264 578212 373316 578264
rect 399024 578212 399076 578264
rect 400864 578212 400916 578264
rect 427360 578212 427412 578264
rect 428556 578212 428608 578264
rect 455328 578212 455380 578264
rect 456064 578212 456116 578264
rect 483204 578212 483256 578264
rect 485044 578212 485096 578264
rect 511356 578212 511408 578264
rect 512644 578212 512696 578264
rect 539324 578212 539376 578264
rect 540244 578212 540296 578264
rect 567200 578212 567252 578264
rect 37924 576104 37976 576156
rect 545764 576104 545816 576156
rect 35624 575424 35676 575476
rect 36728 575424 36780 575476
rect 147680 562300 147732 562352
rect 148416 562300 148468 562352
rect 259736 562300 259788 562352
rect 260196 562300 260248 562352
rect 455696 562300 455748 562352
rect 456156 562300 456208 562352
rect 287704 558832 287756 558884
rect 295708 558832 295760 558884
rect 316776 558832 316828 558884
rect 323676 558832 323728 558884
rect 63592 558288 63644 558340
rect 64328 558288 64380 558340
rect 232688 558152 232740 558204
rect 239772 558152 239824 558204
rect 428648 558152 428700 558204
rect 435732 558152 435784 558204
rect 483664 558152 483716 558204
rect 491668 558152 491720 558204
rect 512736 557608 512788 557660
rect 519636 557608 519688 557660
rect 13728 557472 13780 557524
rect 66260 557472 66312 557524
rect 97908 557472 97960 557524
rect 149060 557472 149112 557524
rect 154488 557472 154540 557524
rect 205640 557472 205692 557524
rect 209688 557472 209740 557524
rect 262220 557472 262272 557524
rect 266268 557472 266320 557524
rect 317420 557472 317472 557524
rect 322848 557472 322900 557524
rect 374000 557472 374052 557524
rect 405648 557472 405700 557524
rect 458180 557472 458232 557524
rect 489828 557472 489880 557524
rect 542360 557472 542412 557524
rect 35624 557404 35676 557456
rect 36912 557404 36964 557456
rect 42708 557404 42760 557456
rect 93860 557404 93912 557456
rect 126888 557404 126940 557456
rect 178040 557404 178092 557456
rect 182088 557404 182140 557456
rect 233240 557404 233292 557456
rect 238668 557404 238720 557456
rect 289820 557404 289872 557456
rect 293868 557404 293920 557456
rect 70308 557336 70360 557388
rect 121460 557336 121512 557388
rect 343548 557404 343600 557456
rect 345664 557404 345716 557456
rect 350448 557404 350500 557456
rect 401600 557404 401652 557456
rect 434628 557404 434680 557456
rect 485780 557404 485832 557456
rect 518808 557404 518860 557456
rect 569960 557404 570012 557456
rect 345020 557336 345072 557388
rect 378048 557336 378100 557388
rect 429200 557336 429252 557388
rect 462228 557336 462280 557388
rect 513380 557336 513432 557388
rect 42892 554684 42944 554736
rect 15200 554616 15252 554668
rect 43996 554616 44048 554668
rect 72056 554684 72108 554736
rect 99472 554684 99524 554736
rect 71872 554616 71924 554668
rect 100024 554616 100076 554668
rect 127072 554684 127124 554736
rect 127992 554616 128044 554668
rect 183652 554684 183704 554736
rect 156052 554616 156104 554668
rect 165988 554616 166040 554668
rect 177304 554616 177356 554668
rect 178684 554616 178736 554668
rect 184020 554616 184072 554668
rect 374644 554684 374696 554736
rect 379704 554684 379756 554736
rect 539324 554684 539376 554736
rect 543004 554684 543056 554736
rect 211712 554616 211764 554668
rect 222016 554616 222068 554668
rect 232596 554616 232648 554668
rect 249708 554616 249760 554668
rect 260104 554616 260156 554668
rect 261484 554616 261536 554668
rect 567200 554616 567252 554668
rect 25688 554548 25740 554600
rect 37004 554548 37056 554600
rect 53656 554548 53708 554600
rect 69664 554548 69716 554600
rect 81992 554548 82044 554600
rect 94504 554548 94556 554600
rect 109684 554548 109736 554600
rect 120724 554548 120776 554600
rect 137652 554548 137704 554600
rect 148324 554548 148376 554600
rect 193680 554548 193732 554600
rect 204904 554548 204956 554600
rect 238852 554548 238904 554600
rect 268016 554548 268068 554600
rect 277676 554548 277728 554600
rect 289084 554548 289136 554600
rect 306012 554548 306064 554600
rect 316684 554548 316736 554600
rect 323032 554548 323084 554600
rect 352012 554548 352064 554600
rect 361672 554548 361724 554600
rect 373264 554548 373316 554600
rect 379612 554548 379664 554600
rect 408040 554548 408092 554600
rect 417700 554548 417752 554600
rect 428556 554548 428608 554600
rect 434812 554548 434864 554600
rect 463700 554548 463752 554600
rect 474004 554548 474056 554600
rect 485044 554548 485096 554600
rect 501696 554548 501748 554600
rect 512644 554548 512696 554600
rect 518992 554548 519044 554600
rect 547880 554548 547932 554600
rect 333704 554480 333756 554532
rect 344284 554480 344336 554532
rect 390008 554480 390060 554532
rect 400864 554480 400916 554532
rect 445668 554480 445720 554532
rect 456064 554480 456116 554532
rect 529664 554480 529716 554532
rect 540244 554480 540296 554532
rect 36820 554412 36872 554464
rect 557540 554412 557592 554464
rect 16028 551284 16080 551336
rect 547880 551284 547932 551336
rect 25688 550876 25740 550928
rect 261484 550876 261536 550928
rect 148324 550808 148376 550860
rect 165712 550808 165764 550860
rect 175464 550808 175516 550860
rect 193680 550808 193732 550860
rect 203524 550808 203576 550860
rect 221372 550808 221424 550860
rect 296352 550808 296404 550860
rect 316776 550808 316828 550860
rect 408040 550808 408092 550860
rect 428648 550808 428700 550860
rect 492036 550808 492088 550860
rect 512736 550808 512788 550860
rect 36820 550740 36872 550792
rect 53656 550740 53708 550792
rect 64328 550740 64380 550792
rect 81440 550740 81492 550792
rect 91468 550740 91520 550792
rect 109684 550740 109736 550792
rect 119436 550740 119488 550792
rect 137652 550740 137704 550792
rect 156328 550740 156380 550792
rect 178684 550740 178736 550792
rect 232504 550740 232556 550792
rect 249708 550740 249760 550792
rect 260104 550740 260156 550792
rect 277676 550740 277728 550792
rect 287520 550740 287572 550792
rect 305368 550740 305420 550792
rect 345664 550740 345716 550792
rect 361672 550740 361724 550792
rect 371516 550740 371568 550792
rect 389364 550740 389416 550792
rect 399484 550740 399536 550792
rect 417700 550740 417752 550792
rect 456156 550740 456208 550792
rect 473360 550740 473412 550792
rect 483480 550740 483532 550792
rect 501696 550740 501748 550792
rect 37004 550672 37056 550724
rect 63316 550672 63368 550724
rect 66904 550672 66956 550724
rect 91100 550672 91152 550724
rect 94504 550672 94556 550724
rect 119344 550672 119396 550724
rect 120724 550672 120776 550724
rect 147312 550672 147364 550724
rect 148416 550672 148468 550724
rect 175372 550672 175424 550724
rect 177304 550672 177356 550724
rect 203340 550672 203392 550724
rect 204904 550672 204956 550724
rect 231032 550672 231084 550724
rect 232596 550672 232648 550724
rect 259368 550672 259420 550724
rect 268016 550672 268068 550724
rect 287704 550672 287756 550724
rect 315488 550672 315540 550724
rect 333704 550672 333756 550724
rect 352012 550672 352064 550724
rect 374644 550672 374696 550724
rect 428464 550672 428516 550724
rect 445668 550672 445720 550724
rect 464344 550672 464396 550724
rect 483664 550672 483716 550724
rect 511448 550672 511500 550724
rect 529664 550672 529716 550724
rect 543004 550672 543056 550724
rect 557540 550672 557592 550724
rect 212356 550604 212408 550656
rect 232688 550604 232740 550656
rect 260196 550604 260248 550656
rect 287336 550604 287388 550656
rect 289084 550604 289136 550656
rect 315028 550604 315080 550656
rect 316684 550604 316736 550656
rect 343364 550604 343416 550656
rect 344284 550604 344336 550656
rect 371332 550604 371384 550656
rect 373264 550604 373316 550656
rect 399024 550604 399076 550656
rect 400864 550604 400916 550656
rect 427360 550604 427412 550656
rect 428556 550604 428608 550656
rect 455328 550604 455380 550656
rect 456064 550604 456116 550656
rect 483020 550604 483072 550656
rect 485044 550604 485096 550656
rect 511356 550604 511408 550656
rect 512644 550604 512696 550656
rect 539324 550604 539376 550656
rect 540244 550604 540296 550656
rect 567200 550604 567252 550656
rect 37924 548496 37976 548548
rect 545764 548496 545816 548548
rect 35624 547884 35676 547936
rect 36912 547884 36964 547936
rect 63592 533604 63644 533656
rect 64328 533604 64380 533656
rect 455696 533604 455748 533656
rect 456156 533604 456208 533656
rect 316776 530680 316828 530732
rect 323676 530680 323728 530732
rect 428648 530544 428700 530596
rect 435732 530544 435784 530596
rect 287704 530272 287756 530324
rect 295708 530272 295760 530324
rect 232688 530204 232740 530256
rect 239772 530204 239824 530256
rect 512736 530204 512788 530256
rect 519636 530204 519688 530256
rect 483664 530136 483716 530188
rect 491668 530136 491720 530188
rect 13728 529864 13780 529916
rect 66260 529864 66312 529916
rect 97908 529864 97960 529916
rect 149060 529864 149112 529916
rect 154488 529864 154540 529916
rect 205640 529864 205692 529916
rect 209688 529864 209740 529916
rect 262220 529864 262272 529916
rect 266268 529864 266320 529916
rect 317420 529864 317472 529916
rect 322848 529864 322900 529916
rect 374000 529864 374052 529916
rect 405648 529864 405700 529916
rect 458180 529864 458232 529916
rect 489828 529864 489880 529916
rect 542360 529864 542412 529916
rect 35624 529796 35676 529848
rect 36820 529796 36872 529848
rect 42708 529796 42760 529848
rect 93860 529796 93912 529848
rect 126888 529796 126940 529848
rect 178040 529796 178092 529848
rect 182088 529796 182140 529848
rect 233240 529796 233292 529848
rect 238668 529796 238720 529848
rect 289820 529796 289872 529848
rect 293868 529796 293920 529848
rect 70308 529728 70360 529780
rect 121460 529728 121512 529780
rect 343548 529796 343600 529848
rect 345664 529796 345716 529848
rect 350448 529796 350500 529848
rect 401600 529796 401652 529848
rect 434628 529796 434680 529848
rect 485780 529796 485832 529848
rect 518808 529796 518860 529848
rect 569960 529796 570012 529848
rect 345020 529728 345072 529780
rect 378048 529728 378100 529780
rect 429200 529728 429252 529780
rect 462228 529728 462280 529780
rect 513380 529728 513432 529780
rect 178684 527076 178736 527128
rect 184020 527076 184072 527128
rect 374644 527076 374696 527128
rect 379704 527076 379756 527128
rect 539324 527076 539376 527128
rect 543004 527076 543056 527128
rect 15200 527008 15252 527060
rect 43996 527008 44048 527060
rect 71044 527008 71096 527060
rect 567200 527008 567252 527060
rect 25688 526940 25740 526992
rect 37004 526940 37056 526992
rect 53656 526940 53708 526992
rect 66904 526940 66956 526992
rect 71872 526940 71924 526992
rect 100024 526940 100076 526992
rect 42892 526872 42944 526924
rect 71964 526872 72016 526924
rect 81992 526872 82044 526924
rect 94504 526872 94556 526924
rect 99472 526872 99524 526924
rect 127992 526940 128044 526992
rect 109684 526872 109736 526924
rect 120724 526872 120776 526924
rect 127072 526872 127124 526924
rect 155960 526940 156012 526992
rect 165988 526940 166040 526992
rect 177304 526940 177356 526992
rect 183652 526940 183704 526992
rect 211712 526940 211764 526992
rect 221924 526940 221976 526992
rect 232596 526940 232648 526992
rect 238852 526940 238904 526992
rect 268016 526940 268068 526992
rect 277676 526940 277728 526992
rect 289084 526940 289136 526992
rect 306012 526940 306064 526992
rect 316684 526940 316736 526992
rect 323032 526940 323084 526992
rect 352012 526940 352064 526992
rect 361672 526940 361724 526992
rect 373264 526940 373316 526992
rect 379612 526940 379664 526992
rect 408040 526940 408092 526992
rect 417700 526940 417752 526992
rect 428556 526940 428608 526992
rect 434812 526940 434864 526992
rect 463792 526940 463844 526992
rect 474004 526940 474056 526992
rect 485044 526940 485096 526992
rect 501696 526940 501748 526992
rect 512644 526940 512696 526992
rect 518992 526940 519044 526992
rect 547880 526940 547932 526992
rect 137652 526872 137704 526924
rect 148416 526872 148468 526924
rect 193680 526872 193732 526924
rect 204904 526872 204956 526924
rect 249708 526872 249760 526924
rect 260196 526872 260248 526924
rect 333704 526872 333756 526924
rect 344284 526872 344336 526924
rect 390008 526872 390060 526924
rect 400864 526872 400916 526924
rect 445668 526872 445720 526924
rect 456064 526872 456116 526924
rect 529664 526872 529716 526924
rect 540244 526872 540296 526924
rect 36728 526804 36780 526856
rect 557540 526804 557592 526856
rect 16028 523676 16080 523728
rect 547880 523676 547932 523728
rect 25688 523200 25740 523252
rect 71044 523200 71096 523252
rect 212356 523200 212408 523252
rect 232688 523200 232740 523252
rect 296352 523200 296404 523252
rect 316776 523200 316828 523252
rect 408040 523200 408092 523252
rect 428648 523200 428700 523252
rect 492036 523200 492088 523252
rect 512736 523200 512788 523252
rect 36728 523132 36780 523184
rect 53656 523132 53708 523184
rect 148416 523132 148468 523184
rect 165712 523132 165764 523184
rect 175464 523132 175516 523184
rect 193680 523132 193732 523184
rect 203524 523132 203576 523184
rect 221372 523132 221424 523184
rect 260196 523132 260248 523184
rect 277676 523132 277728 523184
rect 287520 523132 287572 523184
rect 305368 523132 305420 523184
rect 345664 523132 345716 523184
rect 361672 523132 361724 523184
rect 371516 523132 371568 523184
rect 389364 523132 389416 523184
rect 399484 523132 399536 523184
rect 417700 523132 417752 523184
rect 456156 523132 456208 523184
rect 473360 523132 473412 523184
rect 483480 523132 483532 523184
rect 501696 523132 501748 523184
rect 37004 523064 37056 523116
rect 63316 523064 63368 523116
rect 64328 523064 64380 523116
rect 81440 523064 81492 523116
rect 91468 523064 91520 523116
rect 109684 523064 109736 523116
rect 119436 523064 119488 523116
rect 137652 523064 137704 523116
rect 156328 523064 156380 523116
rect 178684 523064 178736 523116
rect 232504 523064 232556 523116
rect 249708 523064 249760 523116
rect 268016 523064 268068 523116
rect 287704 523064 287756 523116
rect 315488 523064 315540 523116
rect 333704 523064 333756 523116
rect 352012 523064 352064 523116
rect 374644 523064 374696 523116
rect 428556 523064 428608 523116
rect 445668 523064 445720 523116
rect 464344 523064 464396 523116
rect 483664 523064 483716 523116
rect 511448 523064 511500 523116
rect 529664 523064 529716 523116
rect 543004 523064 543056 523116
rect 557540 523064 557592 523116
rect 69664 522996 69716 523048
rect 91100 522996 91152 523048
rect 94504 522996 94556 523048
rect 119344 522996 119396 523048
rect 120724 522996 120776 523048
rect 147312 522996 147364 523048
rect 148324 522996 148376 523048
rect 175372 522996 175424 523048
rect 177304 522996 177356 523048
rect 203340 522996 203392 523048
rect 204904 522996 204956 523048
rect 231032 522996 231084 523048
rect 232596 522996 232648 523048
rect 259368 522996 259420 523048
rect 260104 522996 260156 523048
rect 287336 522996 287388 523048
rect 289084 522996 289136 523048
rect 315028 522996 315080 523048
rect 316684 522996 316736 523048
rect 343364 522996 343416 523048
rect 344284 522996 344336 523048
rect 371332 522996 371384 523048
rect 373264 522996 373316 523048
rect 399024 522996 399076 523048
rect 400864 522996 400916 523048
rect 427360 522996 427412 523048
rect 428464 522996 428516 523048
rect 455328 522996 455380 523048
rect 456064 522996 456116 523048
rect 483020 522996 483072 523048
rect 485044 522996 485096 523048
rect 511356 522996 511408 523048
rect 512644 522996 512696 523048
rect 539324 522996 539376 523048
rect 540244 522996 540296 523048
rect 567200 522996 567252 523048
rect 37924 522248 37976 522300
rect 545764 522248 545816 522300
rect 35624 521704 35676 521756
rect 36820 521704 36872 521756
rect 42708 520344 42760 520396
rect 93860 520344 93912 520396
rect 155868 520344 155920 520396
rect 205640 520344 205692 520396
rect 238668 520344 238720 520396
rect 289820 520344 289872 520396
rect 322848 520344 322900 520396
rect 374000 520344 374052 520396
rect 434628 520344 434680 520396
rect 485780 520344 485832 520396
rect 13728 520276 13780 520328
rect 66260 520276 66312 520328
rect 70308 520276 70360 520328
rect 121460 520276 121512 520328
rect 126888 520276 126940 520328
rect 178040 520276 178092 520328
rect 209688 520276 209740 520328
rect 262220 520276 262272 520328
rect 293868 520276 293920 520328
rect 345020 520276 345072 520328
rect 350448 520276 350500 520328
rect 401600 520276 401652 520328
rect 407856 520276 407908 520328
rect 458180 520276 458232 520328
rect 518808 520276 518860 520328
rect 569960 520276 570012 520328
rect 154488 518848 154540 518900
rect 155868 518848 155920 518900
rect 540888 509192 540940 509244
rect 542360 509192 542412 509244
rect 63592 505588 63644 505640
rect 64328 505588 64380 505640
rect 147680 505588 147732 505640
rect 148416 505588 148468 505640
rect 259736 505588 259788 505640
rect 260196 505588 260248 505640
rect 455696 505588 455748 505640
rect 456156 505588 456208 505640
rect 287704 504568 287756 504620
rect 295708 504568 295760 504620
rect 428648 504364 428700 504416
rect 435732 504364 435784 504416
rect 483664 504296 483716 504348
rect 491668 504296 491720 504348
rect 512736 504296 512788 504348
rect 519636 504296 519688 504348
rect 232688 504228 232740 504280
rect 239772 504228 239824 504280
rect 316776 503752 316828 503804
rect 323676 503752 323728 503804
rect 97908 503616 97960 503668
rect 149060 503616 149112 503668
rect 182088 503616 182140 503668
rect 233240 503616 233292 503668
rect 266268 503616 266320 503668
rect 317420 503616 317472 503668
rect 378048 503616 378100 503668
rect 429200 503616 429252 503668
rect 489828 503616 489880 503668
rect 542360 503616 542412 503668
rect 427728 503548 427780 503600
rect 428556 503548 428608 503600
rect 462228 503548 462280 503600
rect 513380 503548 513432 503600
rect 35624 502256 35676 502308
rect 36728 502256 36780 502308
rect 42892 500896 42944 500948
rect 15200 500828 15252 500880
rect 43996 500828 44048 500880
rect 72056 500896 72108 500948
rect 99472 500896 99524 500948
rect 71872 500828 71924 500880
rect 100024 500828 100076 500880
rect 127072 500896 127124 500948
rect 127992 500828 128044 500880
rect 183652 500896 183704 500948
rect 156052 500828 156104 500880
rect 165988 500828 166040 500880
rect 177304 500828 177356 500880
rect 178684 500828 178736 500880
rect 184020 500828 184072 500880
rect 343364 500896 343416 500948
rect 345664 500896 345716 500948
rect 374644 500896 374696 500948
rect 379704 500896 379756 500948
rect 539324 500896 539376 500948
rect 543004 500896 543056 500948
rect 211712 500828 211764 500880
rect 222016 500828 222068 500880
rect 232596 500828 232648 500880
rect 249708 500828 249760 500880
rect 260104 500828 260156 500880
rect 261484 500828 261536 500880
rect 567200 500828 567252 500880
rect 25688 500760 25740 500812
rect 37004 500760 37056 500812
rect 53656 500760 53708 500812
rect 69664 500760 69716 500812
rect 81992 500760 82044 500812
rect 94504 500760 94556 500812
rect 109684 500760 109736 500812
rect 120724 500760 120776 500812
rect 137652 500760 137704 500812
rect 148324 500760 148376 500812
rect 193680 500760 193732 500812
rect 204904 500760 204956 500812
rect 238852 500760 238904 500812
rect 268016 500760 268068 500812
rect 277676 500760 277728 500812
rect 289084 500760 289136 500812
rect 306012 500760 306064 500812
rect 316684 500760 316736 500812
rect 323032 500760 323084 500812
rect 352012 500760 352064 500812
rect 361672 500760 361724 500812
rect 373264 500760 373316 500812
rect 379612 500760 379664 500812
rect 408040 500760 408092 500812
rect 417700 500760 417752 500812
rect 428464 500760 428516 500812
rect 434812 500760 434864 500812
rect 463700 500760 463752 500812
rect 474004 500760 474056 500812
rect 485044 500760 485096 500812
rect 501696 500760 501748 500812
rect 512644 500760 512696 500812
rect 518992 500760 519044 500812
rect 547880 500760 547932 500812
rect 333704 500692 333756 500744
rect 344284 500692 344336 500744
rect 390008 500692 390060 500744
rect 400864 500692 400916 500744
rect 445668 500692 445720 500744
rect 456064 500692 456116 500744
rect 529664 500692 529716 500744
rect 540244 500692 540296 500744
rect 36912 500624 36964 500676
rect 557540 500624 557592 500676
rect 16028 497428 16080 497480
rect 547880 497428 547932 497480
rect 25688 497088 25740 497140
rect 261484 497088 261536 497140
rect 148416 497020 148468 497072
rect 165712 497020 165764 497072
rect 175464 497020 175516 497072
rect 193680 497020 193732 497072
rect 203524 497020 203576 497072
rect 221372 497020 221424 497072
rect 408040 497020 408092 497072
rect 428648 497020 428700 497072
rect 492036 497020 492088 497072
rect 512736 497020 512788 497072
rect 37004 496952 37056 497004
rect 53656 496952 53708 497004
rect 64328 496952 64380 497004
rect 81440 496952 81492 497004
rect 91468 496952 91520 497004
rect 109684 496952 109736 497004
rect 119436 496952 119488 497004
rect 137652 496952 137704 497004
rect 156328 496952 156380 497004
rect 178684 496952 178736 497004
rect 232504 496952 232556 497004
rect 249708 496952 249760 497004
rect 260104 496952 260156 497004
rect 277676 496952 277728 497004
rect 287520 496952 287572 497004
rect 305368 496952 305420 497004
rect 315488 496952 315540 497004
rect 333704 496952 333756 497004
rect 345664 496952 345716 497004
rect 361672 496952 361724 497004
rect 371516 496952 371568 497004
rect 389364 496952 389416 497004
rect 399484 496952 399536 497004
rect 417700 496952 417752 497004
rect 456156 496952 456208 497004
rect 473360 496952 473412 497004
rect 483480 496952 483532 497004
rect 501696 496952 501748 497004
rect 36912 496884 36964 496936
rect 63316 496884 63368 496936
rect 66904 496884 66956 496936
rect 91100 496884 91152 496936
rect 94504 496884 94556 496936
rect 119344 496884 119396 496936
rect 120724 496884 120776 496936
rect 147312 496884 147364 496936
rect 148324 496884 148376 496936
rect 175372 496884 175424 496936
rect 177304 496884 177356 496936
rect 203340 496884 203392 496936
rect 204904 496884 204956 496936
rect 231032 496884 231084 496936
rect 232596 496884 232648 496936
rect 259368 496884 259420 496936
rect 268016 496884 268068 496936
rect 287704 496884 287756 496936
rect 296352 496884 296404 496936
rect 316776 496884 316828 496936
rect 352012 496884 352064 496936
rect 374644 496884 374696 496936
rect 428556 496884 428608 496936
rect 445668 496884 445720 496936
rect 464344 496884 464396 496936
rect 483664 496884 483716 496936
rect 511448 496884 511500 496936
rect 529664 496884 529716 496936
rect 543004 496884 543056 496936
rect 557540 496884 557592 496936
rect 212356 496816 212408 496868
rect 232688 496816 232740 496868
rect 260196 496816 260248 496868
rect 287336 496816 287388 496868
rect 289084 496816 289136 496868
rect 315028 496816 315080 496868
rect 316684 496816 316736 496868
rect 343364 496816 343416 496868
rect 344284 496816 344336 496868
rect 371332 496816 371384 496868
rect 373264 496816 373316 496868
rect 399024 496816 399076 496868
rect 400864 496816 400916 496868
rect 427360 496816 427412 496868
rect 428464 496816 428516 496868
rect 455328 496816 455380 496868
rect 456064 496816 456116 496868
rect 483020 496816 483072 496868
rect 485044 496816 485096 496868
rect 511356 496816 511408 496868
rect 512644 496816 512696 496868
rect 539324 496816 539376 496868
rect 540244 496816 540296 496868
rect 567200 496816 567252 496868
rect 37924 494708 37976 494760
rect 545764 494708 545816 494760
rect 35624 494028 35676 494080
rect 36728 494028 36780 494080
rect 63592 477640 63644 477692
rect 64328 477640 64380 477692
rect 147680 477640 147732 477692
rect 148416 477640 148468 477692
rect 455696 477640 455748 477692
rect 456156 477640 456208 477692
rect 512736 476960 512788 477012
rect 519636 476960 519688 477012
rect 428648 476756 428700 476808
rect 435732 476756 435784 476808
rect 232688 476552 232740 476604
rect 239772 476552 239824 476604
rect 287704 476416 287756 476468
rect 295708 476416 295760 476468
rect 316776 476416 316828 476468
rect 323676 476416 323728 476468
rect 483664 476280 483716 476332
rect 491668 476280 491720 476332
rect 13728 476008 13780 476060
rect 66260 476008 66312 476060
rect 70308 476008 70360 476060
rect 121460 476008 121512 476060
rect 126888 476008 126940 476060
rect 178040 476008 178092 476060
rect 209688 476008 209740 476060
rect 262220 476008 262272 476060
rect 266268 476008 266320 476060
rect 317420 476008 317472 476060
rect 322848 476008 322900 476060
rect 374000 476008 374052 476060
rect 405648 476008 405700 476060
rect 458180 476008 458232 476060
rect 489828 476008 489880 476060
rect 542360 476008 542412 476060
rect 35624 475940 35676 475992
rect 37004 475940 37056 475992
rect 42708 475940 42760 475992
rect 93860 475940 93912 475992
rect 97908 475940 97960 475992
rect 149060 475940 149112 475992
rect 154488 475940 154540 475992
rect 205640 475940 205692 475992
rect 238668 475940 238720 475992
rect 289820 475940 289872 475992
rect 293868 475940 293920 475992
rect 345020 475940 345072 475992
rect 350448 475940 350500 475992
rect 401600 475940 401652 475992
rect 427728 475940 427780 475992
rect 428556 475940 428608 475992
rect 434628 475940 434680 475992
rect 485780 475940 485832 475992
rect 518808 475940 518860 475992
rect 569960 475940 570012 475992
rect 182088 475872 182140 475924
rect 233240 475872 233292 475924
rect 343548 475872 343600 475924
rect 345664 475872 345716 475924
rect 378048 475872 378100 475924
rect 429200 475872 429252 475924
rect 462228 475872 462280 475924
rect 513380 475872 513432 475924
rect 539508 475872 539560 475924
rect 543004 475872 543056 475924
rect 178684 473288 178736 473340
rect 184020 473288 184072 473340
rect 374644 473288 374696 473340
rect 379704 473288 379756 473340
rect 15200 473220 15252 473272
rect 43996 473220 44048 473272
rect 71044 473220 71096 473272
rect 567200 473220 567252 473272
rect 25688 473152 25740 473204
rect 36912 473152 36964 473204
rect 53656 473152 53708 473204
rect 66904 473152 66956 473204
rect 71872 473152 71924 473204
rect 100024 473152 100076 473204
rect 42892 473084 42944 473136
rect 72056 473084 72108 473136
rect 81992 473084 82044 473136
rect 94504 473084 94556 473136
rect 99472 473084 99524 473136
rect 127992 473152 128044 473204
rect 109684 473084 109736 473136
rect 120724 473084 120776 473136
rect 127072 473084 127124 473136
rect 156052 473152 156104 473204
rect 165988 473152 166040 473204
rect 177304 473152 177356 473204
rect 183652 473152 183704 473204
rect 211712 473152 211764 473204
rect 222016 473152 222068 473204
rect 232596 473152 232648 473204
rect 238852 473152 238904 473204
rect 268016 473152 268068 473204
rect 277676 473152 277728 473204
rect 289084 473152 289136 473204
rect 306012 473152 306064 473204
rect 316684 473152 316736 473204
rect 323032 473152 323084 473204
rect 352012 473152 352064 473204
rect 361672 473152 361724 473204
rect 373264 473152 373316 473204
rect 379612 473152 379664 473204
rect 408040 473152 408092 473204
rect 417700 473152 417752 473204
rect 428464 473152 428516 473204
rect 434812 473152 434864 473204
rect 463700 473152 463752 473204
rect 474004 473152 474056 473204
rect 485044 473152 485096 473204
rect 501696 473152 501748 473204
rect 512644 473152 512696 473204
rect 518992 473152 519044 473204
rect 547880 473152 547932 473204
rect 137652 473084 137704 473136
rect 148324 473084 148376 473136
rect 193680 473084 193732 473136
rect 204904 473084 204956 473136
rect 249708 473084 249760 473136
rect 260196 473084 260248 473136
rect 333704 473084 333756 473136
rect 344284 473084 344336 473136
rect 390008 473084 390060 473136
rect 400864 473084 400916 473136
rect 445668 473084 445720 473136
rect 456064 473084 456116 473136
rect 529664 473084 529716 473136
rect 540244 473084 540296 473136
rect 36820 473016 36872 473068
rect 557540 473016 557592 473068
rect 15292 469820 15344 469872
rect 547880 469820 547932 469872
rect 25688 469412 25740 469464
rect 71044 469412 71096 469464
rect 296352 469412 296404 469464
rect 316776 469412 316828 469464
rect 408040 469412 408092 469464
rect 428648 469412 428700 469464
rect 37004 469344 37056 469396
rect 53656 469344 53708 469396
rect 148416 469344 148468 469396
rect 165712 469344 165764 469396
rect 175464 469344 175516 469396
rect 193680 469344 193732 469396
rect 203524 469344 203576 469396
rect 221372 469344 221424 469396
rect 232504 469344 232556 469396
rect 249708 469344 249760 469396
rect 260104 469344 260156 469396
rect 277676 469344 277728 469396
rect 287520 469344 287572 469396
rect 305368 469344 305420 469396
rect 345664 469344 345716 469396
rect 361672 469344 361724 469396
rect 371516 469344 371568 469396
rect 389364 469344 389416 469396
rect 399484 469344 399536 469396
rect 417700 469344 417752 469396
rect 456156 469344 456208 469396
rect 473360 469344 473412 469396
rect 483480 469344 483532 469396
rect 501696 469344 501748 469396
rect 511448 469344 511500 469396
rect 529664 469344 529716 469396
rect 36912 469276 36964 469328
rect 63316 469276 63368 469328
rect 64328 469276 64380 469328
rect 81440 469276 81492 469328
rect 91468 469276 91520 469328
rect 109684 469276 109736 469328
rect 119436 469276 119488 469328
rect 137652 469276 137704 469328
rect 156328 469276 156380 469328
rect 178684 469276 178736 469328
rect 212356 469276 212408 469328
rect 232688 469276 232740 469328
rect 268016 469276 268068 469328
rect 287704 469276 287756 469328
rect 315488 469276 315540 469328
rect 333704 469276 333756 469328
rect 352012 469276 352064 469328
rect 374644 469276 374696 469328
rect 428464 469276 428516 469328
rect 445668 469276 445720 469328
rect 464344 469276 464396 469328
rect 483664 469276 483716 469328
rect 492036 469276 492088 469328
rect 512736 469276 512788 469328
rect 543004 469276 543056 469328
rect 557540 469276 557592 469328
rect 69664 469208 69716 469260
rect 91100 469208 91152 469260
rect 94504 469208 94556 469260
rect 119344 469208 119396 469260
rect 120724 469208 120776 469260
rect 147312 469208 147364 469260
rect 148324 469208 148376 469260
rect 175372 469208 175424 469260
rect 177304 469208 177356 469260
rect 203340 469208 203392 469260
rect 204904 469208 204956 469260
rect 231032 469208 231084 469260
rect 232596 469208 232648 469260
rect 259368 469208 259420 469260
rect 260196 469208 260248 469260
rect 287336 469208 287388 469260
rect 289084 469208 289136 469260
rect 315028 469208 315080 469260
rect 316684 469208 316736 469260
rect 343364 469208 343416 469260
rect 344284 469208 344336 469260
rect 371332 469208 371384 469260
rect 373264 469208 373316 469260
rect 399024 469208 399076 469260
rect 400864 469208 400916 469260
rect 427360 469208 427412 469260
rect 428556 469208 428608 469260
rect 455328 469208 455380 469260
rect 456064 469208 456116 469260
rect 483020 469208 483072 469260
rect 485044 469208 485096 469260
rect 511356 469208 511408 469260
rect 512644 469208 512696 469260
rect 539324 469208 539376 469260
rect 540244 469208 540296 469260
rect 567200 469208 567252 469260
rect 37924 468460 37976 468512
rect 545764 468460 545816 468512
rect 182088 466556 182140 466608
rect 233240 466556 233292 466608
rect 350448 466556 350500 466608
rect 401600 466556 401652 466608
rect 462228 466556 462280 466608
rect 513380 466556 513432 466608
rect 35624 466488 35676 466540
rect 36820 466488 36872 466540
rect 42708 466488 42760 466540
rect 93860 466488 93912 466540
rect 97908 466488 97960 466540
rect 149060 466488 149112 466540
rect 154488 466488 154540 466540
rect 205640 466488 205692 466540
rect 238668 466488 238720 466540
rect 289820 466488 289872 466540
rect 293868 466488 293920 466540
rect 345020 466488 345072 466540
rect 378048 466488 378100 466540
rect 429200 466488 429252 466540
rect 434628 466488 434680 466540
rect 485780 466488 485832 466540
rect 518808 466488 518860 466540
rect 569960 466488 570012 466540
rect 13728 466420 13780 466472
rect 66260 466420 66312 466472
rect 70308 466420 70360 466472
rect 121460 466420 121512 466472
rect 126888 466420 126940 466472
rect 178040 466420 178092 466472
rect 209688 466420 209740 466472
rect 262220 466420 262272 466472
rect 266268 466420 266320 466472
rect 317420 466420 317472 466472
rect 322848 466420 322900 466472
rect 374000 466420 374052 466472
rect 405648 466420 405700 466472
rect 458180 466420 458232 466472
rect 489828 466420 489880 466472
rect 542360 466420 542412 466472
rect 428648 450508 428700 450560
rect 435732 450508 435784 450560
rect 512736 450440 512788 450492
rect 519636 450440 519688 450492
rect 483664 450304 483716 450356
rect 491668 450304 491720 450356
rect 232688 449896 232740 449948
rect 239772 449896 239824 449948
rect 287704 449896 287756 449948
rect 295708 449896 295760 449948
rect 316776 449896 316828 449948
rect 323676 449896 323728 449948
rect 63592 449624 63644 449676
rect 64328 449624 64380 449676
rect 455696 449624 455748 449676
rect 456156 449624 456208 449676
rect 35624 448468 35676 448520
rect 37004 448468 37056 448520
rect 147680 448468 147732 448520
rect 148416 448468 148468 448520
rect 343640 448468 343692 448520
rect 345664 448468 345716 448520
rect 539508 448468 539560 448520
rect 543004 448468 543056 448520
rect 42892 445680 42944 445732
rect 15200 445612 15252 445664
rect 43996 445612 44048 445664
rect 72056 445680 72108 445732
rect 99472 445680 99524 445732
rect 71872 445612 71924 445664
rect 100024 445612 100076 445664
rect 127072 445680 127124 445732
rect 127992 445612 128044 445664
rect 183652 445680 183704 445732
rect 156052 445612 156104 445664
rect 165988 445612 166040 445664
rect 177304 445612 177356 445664
rect 178684 445612 178736 445664
rect 184020 445612 184072 445664
rect 374644 445680 374696 445732
rect 379704 445680 379756 445732
rect 211712 445612 211764 445664
rect 222016 445612 222068 445664
rect 232596 445612 232648 445664
rect 249708 445612 249760 445664
rect 260196 445612 260248 445664
rect 261484 445612 261536 445664
rect 567200 445612 567252 445664
rect 25688 445544 25740 445596
rect 36912 445544 36964 445596
rect 53656 445544 53708 445596
rect 69664 445544 69716 445596
rect 81992 445544 82044 445596
rect 94504 445544 94556 445596
rect 109684 445544 109736 445596
rect 120724 445544 120776 445596
rect 137652 445544 137704 445596
rect 148324 445544 148376 445596
rect 193680 445544 193732 445596
rect 204904 445544 204956 445596
rect 238852 445544 238904 445596
rect 268016 445544 268068 445596
rect 277676 445544 277728 445596
rect 289084 445544 289136 445596
rect 306012 445544 306064 445596
rect 316684 445544 316736 445596
rect 323032 445544 323084 445596
rect 352012 445544 352064 445596
rect 361672 445544 361724 445596
rect 373264 445544 373316 445596
rect 379612 445544 379664 445596
rect 408040 445544 408092 445596
rect 417700 445544 417752 445596
rect 428556 445544 428608 445596
rect 434812 445544 434864 445596
rect 463700 445544 463752 445596
rect 474004 445544 474056 445596
rect 485044 445544 485096 445596
rect 501696 445544 501748 445596
rect 512644 445544 512696 445596
rect 518992 445544 519044 445596
rect 547880 445544 547932 445596
rect 333704 445476 333756 445528
rect 344284 445476 344336 445528
rect 390008 445476 390060 445528
rect 400864 445476 400916 445528
rect 445668 445476 445720 445528
rect 456064 445476 456116 445528
rect 529664 445476 529716 445528
rect 540244 445476 540296 445528
rect 36728 445408 36780 445460
rect 557540 445408 557592 445460
rect 16028 443640 16080 443692
rect 547880 443640 547932 443692
rect 25688 443164 25740 443216
rect 69664 443164 69716 443216
rect 212264 443164 212316 443216
rect 232688 443164 232740 443216
rect 296352 443164 296404 443216
rect 316776 443164 316828 443216
rect 408040 443164 408092 443216
rect 428648 443164 428700 443216
rect 492036 443164 492088 443216
rect 512736 443164 512788 443216
rect 36912 443096 36964 443148
rect 53380 443096 53432 443148
rect 64328 443096 64380 443148
rect 81440 443096 81492 443148
rect 148324 443096 148376 443148
rect 165620 443096 165672 443148
rect 175464 443096 175516 443148
rect 193680 443096 193732 443148
rect 203524 443096 203576 443148
rect 221372 443096 221424 443148
rect 260196 443096 260248 443148
rect 277676 443096 277728 443148
rect 287520 443096 287572 443148
rect 305368 443096 305420 443148
rect 345664 443096 345716 443148
rect 361672 443096 361724 443148
rect 371516 443096 371568 443148
rect 389364 443096 389416 443148
rect 399484 443096 399536 443148
rect 417700 443096 417752 443148
rect 456064 443096 456116 443148
rect 473544 443096 473596 443148
rect 483480 443096 483532 443148
rect 501696 443096 501748 443148
rect 37004 443028 37056 443080
rect 62948 443028 63000 443080
rect 66904 443028 66956 443080
rect 91100 443028 91152 443080
rect 91468 443028 91520 443080
rect 109684 443028 109736 443080
rect 119436 443028 119488 443080
rect 137284 443028 137336 443080
rect 156328 443028 156380 443080
rect 178684 443028 178736 443080
rect 232504 443028 232556 443080
rect 249340 443028 249392 443080
rect 268016 443028 268068 443080
rect 287704 443028 287756 443080
rect 315488 443028 315540 443080
rect 333428 443028 333480 443080
rect 352012 443028 352064 443080
rect 374644 443028 374696 443080
rect 428556 443028 428608 443080
rect 445668 443028 445720 443080
rect 464344 443028 464396 443080
rect 483664 443028 483716 443080
rect 511448 443028 511500 443080
rect 529664 443028 529716 443080
rect 543004 443028 543056 443080
rect 557540 443028 557592 443080
rect 94504 442960 94556 443012
rect 119344 442960 119396 443012
rect 120724 442960 120776 443012
rect 147036 442960 147088 443012
rect 148416 442960 148468 443012
rect 175280 442960 175332 443012
rect 177304 442960 177356 443012
rect 203340 442960 203392 443012
rect 204904 442960 204956 443012
rect 231032 442960 231084 443012
rect 232596 442960 232648 443012
rect 259092 442960 259144 443012
rect 260104 442960 260156 443012
rect 287336 442960 287388 443012
rect 289084 442960 289136 443012
rect 315028 442960 315080 443012
rect 316684 442960 316736 443012
rect 342996 442960 343048 443012
rect 344284 442960 344336 443012
rect 371332 442960 371384 443012
rect 373264 442960 373316 443012
rect 399024 442960 399076 443012
rect 400864 442960 400916 443012
rect 427360 442960 427412 443012
rect 428464 442960 428516 443012
rect 455328 442960 455380 443012
rect 456156 442960 456208 443012
rect 483204 442960 483256 443012
rect 485044 442960 485096 443012
rect 511356 442960 511408 443012
rect 512644 442960 512696 443012
rect 539324 442960 539376 443012
rect 540244 442960 540296 443012
rect 567200 442960 567252 443012
rect 37924 440852 37976 440904
rect 545764 440852 545816 440904
rect 182088 440308 182140 440360
rect 233240 440308 233292 440360
rect 350448 440308 350500 440360
rect 401600 440308 401652 440360
rect 35624 440240 35676 440292
rect 36728 440240 36780 440292
rect 42708 440240 42760 440292
rect 93860 440240 93912 440292
rect 97908 440240 97960 440292
rect 149060 440240 149112 440292
rect 154488 440240 154540 440292
rect 205640 440240 205692 440292
rect 238668 440240 238720 440292
rect 289820 440240 289872 440292
rect 293868 440240 293920 440292
rect 345020 440240 345072 440292
rect 378048 440240 378100 440292
rect 429200 440240 429252 440292
rect 434628 440240 434680 440292
rect 485780 440240 485832 440292
rect 489828 440240 489880 440292
rect 542360 440240 542412 440292
rect 63592 427116 63644 427168
rect 64328 427116 64380 427168
rect 259736 427116 259788 427168
rect 260196 427116 260248 427168
rect 287704 423580 287756 423632
rect 295708 423580 295760 423632
rect 316776 423580 316828 423632
rect 323676 423580 323728 423632
rect 483664 423036 483716 423088
rect 491668 423036 491720 423088
rect 232688 422968 232740 423020
rect 239772 422968 239824 423020
rect 512736 422968 512788 423020
rect 519636 422968 519688 423020
rect 428648 422900 428700 422952
rect 435732 422900 435784 422952
rect 13728 422220 13780 422272
rect 66260 422220 66312 422272
rect 70308 422220 70360 422272
rect 121460 422220 121512 422272
rect 126888 422220 126940 422272
rect 178040 422220 178092 422272
rect 209688 422220 209740 422272
rect 262220 422220 262272 422272
rect 266268 422220 266320 422272
rect 317420 422220 317472 422272
rect 322848 422220 322900 422272
rect 374000 422220 374052 422272
rect 405648 422220 405700 422272
rect 458180 422220 458232 422272
rect 462228 422220 462280 422272
rect 513380 422220 513432 422272
rect 518808 422220 518860 422272
rect 569960 422220 570012 422272
rect 35624 422152 35676 422204
rect 36912 422152 36964 422204
rect 343548 422152 343600 422204
rect 345664 422152 345716 422204
rect 427728 421676 427780 421728
rect 428556 421676 428608 421728
rect 539508 421676 539560 421728
rect 543004 421676 543056 421728
rect 178684 419432 178736 419484
rect 184020 419432 184072 419484
rect 374644 419432 374696 419484
rect 379704 419432 379756 419484
rect 15200 419364 15252 419416
rect 43996 419364 44048 419416
rect 71044 419364 71096 419416
rect 567200 419364 567252 419416
rect 25688 419296 25740 419348
rect 37004 419296 37056 419348
rect 53656 419296 53708 419348
rect 66904 419296 66956 419348
rect 71872 419296 71924 419348
rect 100024 419296 100076 419348
rect 42892 419228 42944 419280
rect 72056 419228 72108 419280
rect 81992 419228 82044 419280
rect 94504 419228 94556 419280
rect 99472 419228 99524 419280
rect 127992 419296 128044 419348
rect 109684 419228 109736 419280
rect 120724 419228 120776 419280
rect 127072 419228 127124 419280
rect 156052 419296 156104 419348
rect 165988 419296 166040 419348
rect 177304 419296 177356 419348
rect 183652 419296 183704 419348
rect 211712 419296 211764 419348
rect 222016 419296 222068 419348
rect 232596 419296 232648 419348
rect 238852 419296 238904 419348
rect 268016 419296 268068 419348
rect 277676 419296 277728 419348
rect 289084 419296 289136 419348
rect 306012 419296 306064 419348
rect 316684 419296 316736 419348
rect 323032 419296 323084 419348
rect 352012 419296 352064 419348
rect 361672 419296 361724 419348
rect 373264 419296 373316 419348
rect 379612 419296 379664 419348
rect 408040 419296 408092 419348
rect 417700 419296 417752 419348
rect 428464 419296 428516 419348
rect 434812 419296 434864 419348
rect 463700 419296 463752 419348
rect 474004 419296 474056 419348
rect 485044 419296 485096 419348
rect 501696 419296 501748 419348
rect 512644 419296 512696 419348
rect 518992 419296 519044 419348
rect 547880 419296 547932 419348
rect 137652 419228 137704 419280
rect 148416 419228 148468 419280
rect 193680 419228 193732 419280
rect 204904 419228 204956 419280
rect 249708 419228 249760 419280
rect 260104 419228 260156 419280
rect 333704 419228 333756 419280
rect 344284 419228 344336 419280
rect 390008 419228 390060 419280
rect 400864 419228 400916 419280
rect 445668 419228 445720 419280
rect 456156 419228 456208 419280
rect 529664 419228 529716 419280
rect 540244 419228 540296 419280
rect 36820 419160 36872 419212
rect 557540 419160 557592 419212
rect 16028 416032 16080 416084
rect 547880 416032 547932 416084
rect 25688 415692 25740 415744
rect 261484 415692 261536 415744
rect 119436 415624 119488 415676
rect 137652 415624 137704 415676
rect 148324 415624 148376 415676
rect 165712 415624 165764 415676
rect 175464 415624 175516 415676
rect 193680 415624 193732 415676
rect 203524 415624 203576 415676
rect 221372 415624 221424 415676
rect 408040 415624 408092 415676
rect 428648 415624 428700 415676
rect 492036 415624 492088 415676
rect 512736 415624 512788 415676
rect 37004 415556 37056 415608
rect 53656 415556 53708 415608
rect 64328 415556 64380 415608
rect 81440 415556 81492 415608
rect 91468 415556 91520 415608
rect 109684 415556 109736 415608
rect 127992 415556 128044 415608
rect 148508 415556 148560 415608
rect 156328 415556 156380 415608
rect 178684 415556 178736 415608
rect 232596 415556 232648 415608
rect 249708 415556 249760 415608
rect 260196 415556 260248 415608
rect 277676 415556 277728 415608
rect 287520 415556 287572 415608
rect 305368 415556 305420 415608
rect 315488 415556 315540 415608
rect 333704 415556 333756 415608
rect 345664 415556 345716 415608
rect 361672 415556 361724 415608
rect 371516 415556 371568 415608
rect 389364 415556 389416 415608
rect 399484 415556 399536 415608
rect 417700 415556 417752 415608
rect 456156 415556 456208 415608
rect 473360 415556 473412 415608
rect 483480 415556 483532 415608
rect 501696 415556 501748 415608
rect 36912 415488 36964 415540
rect 63316 415488 63368 415540
rect 66904 415488 66956 415540
rect 91100 415488 91152 415540
rect 94504 415488 94556 415540
rect 119344 415488 119396 415540
rect 120724 415488 120776 415540
rect 147312 415488 147364 415540
rect 148416 415488 148468 415540
rect 175372 415488 175424 415540
rect 177304 415488 177356 415540
rect 203340 415488 203392 415540
rect 204904 415488 204956 415540
rect 231032 415488 231084 415540
rect 232504 415488 232556 415540
rect 259368 415488 259420 415540
rect 268016 415488 268068 415540
rect 287704 415488 287756 415540
rect 296352 415488 296404 415540
rect 316776 415488 316828 415540
rect 352012 415488 352064 415540
rect 374644 415488 374696 415540
rect 428556 415488 428608 415540
rect 445668 415488 445720 415540
rect 464344 415488 464396 415540
rect 483664 415488 483716 415540
rect 511448 415488 511500 415540
rect 529664 415488 529716 415540
rect 543004 415488 543056 415540
rect 557540 415488 557592 415540
rect 212356 415420 212408 415472
rect 232688 415420 232740 415472
rect 260104 415420 260156 415472
rect 287336 415420 287388 415472
rect 289084 415420 289136 415472
rect 315028 415420 315080 415472
rect 316684 415420 316736 415472
rect 343364 415420 343416 415472
rect 344284 415420 344336 415472
rect 371332 415420 371384 415472
rect 373264 415420 373316 415472
rect 399024 415420 399076 415472
rect 400864 415420 400916 415472
rect 427360 415420 427412 415472
rect 428464 415420 428516 415472
rect 455328 415420 455380 415472
rect 456064 415420 456116 415472
rect 483020 415420 483072 415472
rect 485044 415420 485096 415472
rect 511356 415420 511408 415472
rect 512644 415420 512696 415472
rect 539324 415420 539376 415472
rect 540244 415420 540296 415472
rect 567200 415420 567252 415472
rect 37924 414672 37976 414724
rect 545764 414672 545816 414724
rect 35624 412632 35676 412684
rect 36820 412632 36872 412684
rect 3332 409844 3384 409896
rect 13084 409844 13136 409896
rect 259736 398488 259788 398540
rect 260196 398488 260248 398540
rect 455696 398488 455748 398540
rect 456156 398488 456208 398540
rect 3332 397468 3384 397520
rect 11704 397468 11756 397520
rect 148508 395292 148560 395344
rect 155868 395292 155920 395344
rect 428648 395292 428700 395344
rect 435732 395292 435784 395344
rect 287704 395088 287756 395140
rect 295800 395088 295852 395140
rect 316776 395088 316828 395140
rect 323676 395088 323728 395140
rect 232688 395020 232740 395072
rect 239772 395020 239824 395072
rect 483664 395020 483716 395072
rect 491668 395020 491720 395072
rect 512736 395020 512788 395072
rect 519636 395020 519688 395072
rect 13728 394612 13780 394664
rect 35624 394544 35676 394596
rect 37004 394544 37056 394596
rect 42708 394544 42760 394596
rect 63592 394612 63644 394664
rect 64328 394612 64380 394664
rect 70308 394612 70360 394664
rect 121460 394612 121512 394664
rect 126888 394612 126940 394664
rect 178040 394612 178092 394664
rect 209688 394612 209740 394664
rect 262220 394612 262272 394664
rect 266268 394612 266320 394664
rect 317420 394612 317472 394664
rect 322848 394612 322900 394664
rect 374000 394612 374052 394664
rect 405648 394612 405700 394664
rect 458180 394612 458232 394664
rect 489828 394612 489880 394664
rect 542360 394612 542412 394664
rect 66260 394476 66312 394528
rect 93860 394544 93912 394596
rect 97908 394544 97960 394596
rect 149060 394544 149112 394596
rect 182088 394544 182140 394596
rect 233240 394544 233292 394596
rect 238668 394544 238720 394596
rect 289820 394544 289872 394596
rect 293868 394544 293920 394596
rect 154488 394476 154540 394528
rect 205640 394476 205692 394528
rect 343640 394544 343692 394596
rect 345664 394544 345716 394596
rect 350448 394544 350500 394596
rect 401600 394544 401652 394596
rect 427728 394544 427780 394596
rect 428556 394544 428608 394596
rect 462228 394544 462280 394596
rect 513380 394544 513432 394596
rect 518808 394544 518860 394596
rect 569960 394544 570012 394596
rect 345020 394476 345072 394528
rect 378048 394476 378100 394528
rect 429200 394476 429252 394528
rect 434628 394476 434680 394528
rect 485780 394476 485832 394528
rect 231584 393252 231636 393304
rect 232596 393252 232648 393304
rect 25688 391892 25740 391944
rect 36912 391892 36964 391944
rect 178684 391892 178736 391944
rect 184020 391892 184072 391944
rect 374644 391892 374696 391944
rect 379704 391892 379756 391944
rect 539324 391892 539376 391944
rect 543004 391892 543056 391944
rect 15200 391824 15252 391876
rect 43996 391824 44048 391876
rect 69664 391824 69716 391876
rect 567200 391824 567252 391876
rect 53656 391756 53708 391808
rect 66904 391756 66956 391808
rect 71872 391756 71924 391808
rect 100024 391756 100076 391808
rect 42892 391688 42944 391740
rect 71964 391688 72016 391740
rect 81992 391688 82044 391740
rect 94504 391688 94556 391740
rect 99472 391688 99524 391740
rect 127992 391756 128044 391808
rect 137652 391756 137704 391808
rect 148416 391756 148468 391808
rect 165988 391756 166040 391808
rect 177304 391756 177356 391808
rect 183652 391756 183704 391808
rect 211712 391756 211764 391808
rect 221924 391756 221976 391808
rect 232504 391756 232556 391808
rect 238852 391756 238904 391808
rect 268016 391756 268068 391808
rect 277676 391756 277728 391808
rect 289084 391756 289136 391808
rect 306012 391756 306064 391808
rect 316684 391756 316736 391808
rect 323032 391756 323084 391808
rect 352012 391756 352064 391808
rect 361672 391756 361724 391808
rect 373264 391756 373316 391808
rect 379612 391756 379664 391808
rect 408040 391756 408092 391808
rect 417700 391756 417752 391808
rect 428464 391756 428516 391808
rect 434812 391756 434864 391808
rect 463792 391756 463844 391808
rect 474004 391756 474056 391808
rect 485044 391756 485096 391808
rect 501696 391756 501748 391808
rect 512644 391756 512696 391808
rect 518992 391756 519044 391808
rect 547880 391756 547932 391808
rect 109684 391688 109736 391740
rect 120724 391688 120776 391740
rect 193680 391688 193732 391740
rect 204904 391688 204956 391740
rect 249708 391688 249760 391740
rect 260104 391688 260156 391740
rect 333704 391688 333756 391740
rect 344284 391688 344336 391740
rect 390008 391688 390060 391740
rect 400864 391688 400916 391740
rect 445668 391688 445720 391740
rect 456064 391688 456116 391740
rect 529664 391688 529716 391740
rect 540244 391688 540296 391740
rect 36728 391620 36780 391672
rect 557540 391620 557592 391672
rect 16028 389784 16080 389836
rect 547880 389784 547932 389836
rect 25688 389376 25740 389428
rect 71044 389376 71096 389428
rect 212356 389376 212408 389428
rect 232688 389376 232740 389428
rect 296352 389376 296404 389428
rect 316776 389376 316828 389428
rect 408040 389376 408092 389428
rect 428648 389376 428700 389428
rect 492036 389376 492088 389428
rect 512736 389376 512788 389428
rect 37004 389308 37056 389360
rect 53656 389308 53708 389360
rect 148416 389308 148468 389360
rect 165712 389308 165764 389360
rect 175464 389308 175516 389360
rect 193680 389308 193732 389360
rect 203524 389308 203576 389360
rect 221372 389308 221424 389360
rect 260104 389308 260156 389360
rect 277676 389308 277728 389360
rect 287520 389308 287572 389360
rect 305368 389308 305420 389360
rect 345664 389308 345716 389360
rect 361672 389308 361724 389360
rect 371516 389308 371568 389360
rect 389364 389308 389416 389360
rect 399484 389308 399536 389360
rect 417700 389308 417752 389360
rect 456156 389308 456208 389360
rect 473360 389308 473412 389360
rect 483480 389308 483532 389360
rect 501696 389308 501748 389360
rect 36912 389240 36964 389292
rect 63316 389240 63368 389292
rect 64328 389240 64380 389292
rect 81440 389240 81492 389292
rect 91468 389240 91520 389292
rect 109684 389240 109736 389292
rect 119436 389240 119488 389292
rect 137652 389240 137704 389292
rect 156328 389240 156380 389292
rect 178684 389240 178736 389292
rect 232596 389240 232648 389292
rect 249708 389240 249760 389292
rect 268016 389240 268068 389292
rect 287704 389240 287756 389292
rect 315488 389240 315540 389292
rect 333704 389240 333756 389292
rect 352012 389240 352064 389292
rect 374644 389240 374696 389292
rect 428556 389240 428608 389292
rect 445668 389240 445720 389292
rect 464344 389240 464396 389292
rect 483664 389240 483716 389292
rect 511448 389240 511500 389292
rect 529664 389240 529716 389292
rect 543004 389240 543056 389292
rect 557540 389240 557592 389292
rect 69664 389172 69716 389224
rect 91100 389172 91152 389224
rect 94504 389172 94556 389224
rect 119344 389172 119396 389224
rect 120724 389172 120776 389224
rect 147312 389172 147364 389224
rect 148324 389172 148376 389224
rect 175372 389172 175424 389224
rect 177304 389172 177356 389224
rect 203340 389172 203392 389224
rect 204904 389172 204956 389224
rect 231032 389172 231084 389224
rect 232504 389172 232556 389224
rect 259368 389172 259420 389224
rect 260196 389172 260248 389224
rect 287336 389172 287388 389224
rect 289084 389172 289136 389224
rect 315028 389172 315080 389224
rect 316684 389172 316736 389224
rect 343364 389172 343416 389224
rect 344284 389172 344336 389224
rect 371332 389172 371384 389224
rect 373264 389172 373316 389224
rect 399024 389172 399076 389224
rect 400864 389172 400916 389224
rect 427360 389172 427412 389224
rect 428464 389172 428516 389224
rect 455328 389172 455380 389224
rect 456064 389172 456116 389224
rect 483020 389172 483072 389224
rect 485044 389172 485096 389224
rect 511356 389172 511408 389224
rect 512644 389172 512696 389224
rect 539324 389172 539376 389224
rect 540244 389172 540296 389224
rect 567200 389172 567252 389224
rect 37924 387064 37976 387116
rect 545764 387064 545816 387116
rect 35624 386384 35676 386436
rect 36728 386384 36780 386436
rect 63592 370540 63644 370592
rect 64328 370540 64380 370592
rect 147680 370540 147732 370592
rect 148416 370540 148468 370592
rect 455696 370540 455748 370592
rect 456156 370540 456208 370592
rect 232688 369248 232740 369300
rect 239772 369248 239824 369300
rect 428648 369112 428700 369164
rect 435732 369112 435784 369164
rect 287704 368840 287756 368892
rect 295708 368840 295760 368892
rect 316776 368840 316828 368892
rect 323676 368840 323728 368892
rect 483664 368840 483716 368892
rect 491668 368840 491720 368892
rect 512736 368704 512788 368756
rect 519636 368704 519688 368756
rect 13728 368432 13780 368484
rect 66260 368432 66312 368484
rect 70308 368432 70360 368484
rect 121460 368432 121512 368484
rect 126888 368432 126940 368484
rect 178040 368432 178092 368484
rect 209688 368432 209740 368484
rect 260748 368432 260800 368484
rect 266268 368432 266320 368484
rect 317420 368432 317472 368484
rect 322848 368432 322900 368484
rect 374000 368432 374052 368484
rect 405648 368432 405700 368484
rect 458180 368432 458232 368484
rect 489828 368432 489880 368484
rect 540888 368432 540940 368484
rect 42708 368364 42760 368416
rect 93860 368364 93912 368416
rect 97908 368364 97960 368416
rect 149060 368364 149112 368416
rect 182088 368364 182140 368416
rect 233240 368364 233292 368416
rect 238668 368364 238720 368416
rect 289820 368364 289872 368416
rect 293868 368364 293920 368416
rect 345020 368364 345072 368416
rect 378048 368364 378100 368416
rect 429200 368364 429252 368416
rect 462228 368364 462280 368416
rect 513380 368364 513432 368416
rect 518808 368364 518860 368416
rect 569960 368364 570012 368416
rect 154488 368296 154540 368348
rect 205640 368296 205692 368348
rect 231676 368296 231728 368348
rect 232596 368296 232648 368348
rect 350448 368296 350500 368348
rect 401600 368296 401652 368348
rect 427728 368296 427780 368348
rect 428556 368296 428608 368348
rect 434628 368296 434680 368348
rect 485780 368296 485832 368348
rect 35624 367004 35676 367056
rect 37004 367004 37056 367056
rect 343548 367004 343600 367056
rect 345664 367004 345716 367056
rect 25688 365644 25740 365696
rect 36912 365644 36964 365696
rect 42892 365644 42944 365696
rect 15200 365576 15252 365628
rect 43996 365576 44048 365628
rect 72056 365644 72108 365696
rect 99472 365644 99524 365696
rect 71872 365576 71924 365628
rect 100024 365576 100076 365628
rect 127072 365644 127124 365696
rect 127992 365576 128044 365628
rect 183652 365644 183704 365696
rect 156052 365576 156104 365628
rect 165988 365576 166040 365628
rect 177304 365576 177356 365628
rect 178684 365576 178736 365628
rect 184020 365576 184072 365628
rect 374644 365644 374696 365696
rect 379704 365644 379756 365696
rect 539324 365644 539376 365696
rect 543004 365644 543056 365696
rect 211712 365576 211764 365628
rect 222016 365576 222068 365628
rect 232504 365576 232556 365628
rect 249708 365576 249760 365628
rect 260196 365576 260248 365628
rect 261484 365576 261536 365628
rect 567200 365576 567252 365628
rect 53656 365508 53708 365560
rect 69664 365508 69716 365560
rect 81992 365508 82044 365560
rect 94504 365508 94556 365560
rect 109684 365508 109736 365560
rect 120724 365508 120776 365560
rect 137652 365508 137704 365560
rect 148324 365508 148376 365560
rect 193680 365508 193732 365560
rect 204904 365508 204956 365560
rect 238852 365508 238904 365560
rect 268016 365508 268068 365560
rect 277676 365508 277728 365560
rect 289084 365508 289136 365560
rect 306012 365508 306064 365560
rect 316684 365508 316736 365560
rect 323032 365508 323084 365560
rect 352012 365508 352064 365560
rect 361672 365508 361724 365560
rect 373264 365508 373316 365560
rect 379612 365508 379664 365560
rect 408040 365508 408092 365560
rect 417700 365508 417752 365560
rect 428464 365508 428516 365560
rect 434812 365508 434864 365560
rect 463700 365508 463752 365560
rect 474004 365508 474056 365560
rect 485044 365508 485096 365560
rect 501696 365508 501748 365560
rect 512644 365508 512696 365560
rect 518992 365508 519044 365560
rect 547880 365508 547932 365560
rect 333704 365440 333756 365492
rect 344284 365440 344336 365492
rect 390008 365440 390060 365492
rect 400864 365440 400916 365492
rect 445668 365440 445720 365492
rect 456064 365440 456116 365492
rect 529664 365440 529716 365492
rect 540244 365440 540296 365492
rect 36820 365372 36872 365424
rect 557540 365372 557592 365424
rect 16028 362176 16080 362228
rect 547880 362176 547932 362228
rect 25688 361836 25740 361888
rect 261484 361836 261536 361888
rect 148416 361768 148468 361820
rect 165712 361768 165764 361820
rect 175464 361768 175516 361820
rect 193680 361768 193732 361820
rect 203524 361768 203576 361820
rect 221372 361768 221424 361820
rect 296352 361768 296404 361820
rect 316776 361768 316828 361820
rect 408040 361768 408092 361820
rect 428648 361768 428700 361820
rect 492036 361768 492088 361820
rect 512736 361768 512788 361820
rect 37004 361700 37056 361752
rect 53656 361700 53708 361752
rect 64328 361700 64380 361752
rect 81440 361700 81492 361752
rect 91468 361700 91520 361752
rect 109684 361700 109736 361752
rect 119436 361700 119488 361752
rect 137652 361700 137704 361752
rect 156328 361700 156380 361752
rect 178684 361700 178736 361752
rect 232596 361700 232648 361752
rect 249708 361700 249760 361752
rect 260104 361700 260156 361752
rect 277676 361700 277728 361752
rect 287520 361700 287572 361752
rect 305368 361700 305420 361752
rect 345664 361700 345716 361752
rect 361672 361700 361724 361752
rect 371516 361700 371568 361752
rect 389364 361700 389416 361752
rect 399484 361700 399536 361752
rect 417700 361700 417752 361752
rect 456064 361700 456116 361752
rect 473360 361700 473412 361752
rect 483480 361700 483532 361752
rect 501696 361700 501748 361752
rect 36820 361632 36872 361684
rect 63316 361632 63368 361684
rect 66904 361632 66956 361684
rect 91100 361632 91152 361684
rect 94504 361632 94556 361684
rect 119344 361632 119396 361684
rect 120724 361632 120776 361684
rect 147312 361632 147364 361684
rect 148324 361632 148376 361684
rect 175372 361632 175424 361684
rect 177304 361632 177356 361684
rect 203340 361632 203392 361684
rect 204904 361632 204956 361684
rect 231032 361632 231084 361684
rect 232504 361632 232556 361684
rect 259368 361632 259420 361684
rect 268016 361632 268068 361684
rect 287704 361632 287756 361684
rect 315488 361632 315540 361684
rect 333704 361632 333756 361684
rect 352012 361632 352064 361684
rect 374644 361632 374696 361684
rect 428556 361632 428608 361684
rect 445668 361632 445720 361684
rect 464344 361632 464396 361684
rect 483664 361632 483716 361684
rect 511448 361632 511500 361684
rect 529664 361632 529716 361684
rect 543004 361632 543056 361684
rect 557540 361632 557592 361684
rect 212356 361564 212408 361616
rect 232688 361564 232740 361616
rect 260196 361564 260248 361616
rect 287336 361564 287388 361616
rect 289084 361564 289136 361616
rect 315028 361564 315080 361616
rect 316684 361564 316736 361616
rect 343364 361564 343416 361616
rect 344284 361564 344336 361616
rect 371332 361564 371384 361616
rect 373264 361564 373316 361616
rect 399024 361564 399076 361616
rect 400864 361564 400916 361616
rect 427360 361564 427412 361616
rect 428464 361564 428516 361616
rect 455328 361564 455380 361616
rect 456156 361564 456208 361616
rect 483020 361564 483072 361616
rect 485044 361564 485096 361616
rect 511356 361564 511408 361616
rect 512644 361564 512696 361616
rect 539324 361564 539376 361616
rect 540244 361564 540296 361616
rect 567200 361564 567252 361616
rect 37924 359456 37976 359508
rect 545764 359456 545816 359508
rect 35624 358776 35676 358828
rect 36912 358776 36964 358828
rect 3332 357416 3384 357468
rect 14464 357416 14516 357468
rect 63592 342524 63644 342576
rect 64328 342524 64380 342576
rect 147680 342524 147732 342576
rect 148416 342524 148468 342576
rect 316776 341912 316828 341964
rect 323676 341912 323728 341964
rect 512736 341912 512788 341964
rect 519636 341912 519688 341964
rect 287704 341504 287756 341556
rect 295708 341504 295760 341556
rect 428648 341504 428700 341556
rect 435732 341504 435784 341556
rect 232688 341368 232740 341420
rect 239772 341368 239824 341420
rect 483664 341368 483716 341420
rect 491668 341368 491720 341420
rect 13728 340824 13780 340876
rect 66260 340824 66312 340876
rect 70308 340824 70360 340876
rect 121460 340824 121512 340876
rect 126888 340824 126940 340876
rect 178040 340824 178092 340876
rect 209688 340824 209740 340876
rect 262220 340824 262272 340876
rect 266268 340824 266320 340876
rect 317420 340824 317472 340876
rect 322848 340824 322900 340876
rect 374000 340824 374052 340876
rect 405648 340824 405700 340876
rect 458180 340824 458232 340876
rect 489828 340824 489880 340876
rect 542360 340824 542412 340876
rect 35624 340756 35676 340808
rect 37004 340756 37056 340808
rect 42708 340756 42760 340808
rect 93860 340756 93912 340808
rect 97908 340756 97960 340808
rect 149060 340756 149112 340808
rect 154488 340756 154540 340808
rect 205640 340756 205692 340808
rect 231676 340756 231728 340808
rect 232596 340756 232648 340808
rect 238668 340756 238720 340808
rect 289820 340756 289872 340808
rect 293868 340756 293920 340808
rect 345020 340756 345072 340808
rect 350448 340756 350500 340808
rect 401600 340756 401652 340808
rect 427728 340756 427780 340808
rect 428556 340756 428608 340808
rect 434628 340756 434680 340808
rect 485780 340756 485832 340808
rect 518808 340756 518860 340808
rect 569960 340756 570012 340808
rect 182088 340688 182140 340740
rect 233240 340688 233292 340740
rect 343640 340688 343692 340740
rect 345664 340688 345716 340740
rect 378048 340688 378100 340740
rect 429200 340688 429252 340740
rect 462228 340688 462280 340740
rect 513380 340688 513432 340740
rect 539508 340688 539560 340740
rect 543004 340688 543056 340740
rect 178684 338036 178736 338088
rect 184020 338036 184072 338088
rect 374644 338036 374696 338088
rect 379704 338036 379756 338088
rect 15200 337968 15252 338020
rect 43996 337968 44048 338020
rect 71044 337968 71096 338020
rect 567200 337968 567252 338020
rect 25688 337900 25740 337952
rect 36820 337900 36872 337952
rect 53656 337900 53708 337952
rect 66904 337900 66956 337952
rect 71872 337900 71924 337952
rect 100024 337900 100076 337952
rect 42892 337832 42944 337884
rect 72056 337832 72108 337884
rect 81992 337832 82044 337884
rect 94504 337832 94556 337884
rect 99472 337832 99524 337884
rect 127992 337900 128044 337952
rect 109684 337832 109736 337884
rect 120724 337832 120776 337884
rect 127072 337832 127124 337884
rect 156052 337900 156104 337952
rect 165988 337900 166040 337952
rect 177304 337900 177356 337952
rect 183652 337900 183704 337952
rect 211712 337900 211764 337952
rect 222016 337900 222068 337952
rect 232504 337900 232556 337952
rect 238852 337900 238904 337952
rect 268016 337900 268068 337952
rect 277676 337900 277728 337952
rect 289084 337900 289136 337952
rect 306012 337900 306064 337952
rect 316684 337900 316736 337952
rect 323032 337900 323084 337952
rect 352012 337900 352064 337952
rect 361672 337900 361724 337952
rect 373264 337900 373316 337952
rect 379612 337900 379664 337952
rect 408040 337900 408092 337952
rect 417700 337900 417752 337952
rect 428464 337900 428516 337952
rect 434812 337900 434864 337952
rect 463700 337900 463752 337952
rect 474004 337900 474056 337952
rect 485044 337900 485096 337952
rect 501696 337900 501748 337952
rect 512644 337900 512696 337952
rect 518992 337900 519044 337952
rect 547880 337900 547932 337952
rect 137652 337832 137704 337884
rect 148324 337832 148376 337884
rect 193680 337832 193732 337884
rect 204904 337832 204956 337884
rect 249708 337832 249760 337884
rect 260196 337832 260248 337884
rect 333704 337832 333756 337884
rect 344284 337832 344336 337884
rect 390008 337832 390060 337884
rect 400864 337832 400916 337884
rect 445668 337832 445720 337884
rect 456156 337832 456208 337884
rect 529664 337832 529716 337884
rect 540244 337832 540296 337884
rect 36728 337764 36780 337816
rect 557540 337764 557592 337816
rect 16028 335996 16080 336048
rect 547880 335996 547932 336048
rect 25688 335520 25740 335572
rect 71044 335520 71096 335572
rect 212264 335520 212316 335572
rect 232688 335520 232740 335572
rect 296352 335520 296404 335572
rect 316776 335520 316828 335572
rect 408040 335520 408092 335572
rect 428648 335520 428700 335572
rect 492036 335520 492088 335572
rect 512736 335520 512788 335572
rect 37004 335452 37056 335504
rect 53656 335452 53708 335504
rect 148324 335452 148376 335504
rect 165620 335452 165672 335504
rect 175464 335452 175516 335504
rect 193680 335452 193732 335504
rect 203524 335452 203576 335504
rect 221372 335452 221424 335504
rect 260196 335452 260248 335504
rect 277676 335452 277728 335504
rect 287520 335452 287572 335504
rect 305368 335452 305420 335504
rect 345664 335452 345716 335504
rect 361672 335452 361724 335504
rect 371516 335452 371568 335504
rect 389364 335452 389416 335504
rect 399484 335452 399536 335504
rect 417700 335452 417752 335504
rect 456156 335452 456208 335504
rect 473544 335452 473596 335504
rect 483480 335452 483532 335504
rect 501696 335452 501748 335504
rect 36728 335384 36780 335436
rect 63316 335384 63368 335436
rect 64328 335384 64380 335436
rect 81440 335384 81492 335436
rect 91468 335384 91520 335436
rect 109684 335384 109736 335436
rect 119436 335384 119488 335436
rect 137652 335384 137704 335436
rect 156328 335384 156380 335436
rect 178684 335384 178736 335436
rect 232504 335384 232556 335436
rect 249708 335384 249760 335436
rect 268016 335384 268068 335436
rect 287704 335384 287756 335436
rect 315488 335384 315540 335436
rect 333704 335384 333756 335436
rect 352012 335384 352064 335436
rect 374644 335384 374696 335436
rect 428556 335384 428608 335436
rect 445668 335384 445720 335436
rect 464344 335384 464396 335436
rect 483664 335384 483716 335436
rect 511448 335384 511500 335436
rect 529664 335384 529716 335436
rect 543004 335384 543056 335436
rect 557540 335384 557592 335436
rect 69664 335316 69716 335368
rect 91100 335316 91152 335368
rect 94504 335316 94556 335368
rect 119344 335316 119396 335368
rect 120724 335316 120776 335368
rect 147312 335316 147364 335368
rect 148416 335316 148468 335368
rect 175280 335316 175332 335368
rect 177304 335316 177356 335368
rect 203340 335316 203392 335368
rect 204904 335316 204956 335368
rect 231032 335316 231084 335368
rect 232596 335316 232648 335368
rect 259368 335316 259420 335368
rect 260104 335316 260156 335368
rect 287336 335316 287388 335368
rect 289084 335316 289136 335368
rect 315028 335316 315080 335368
rect 316684 335316 316736 335368
rect 343364 335316 343416 335368
rect 344284 335316 344336 335368
rect 371332 335316 371384 335368
rect 373264 335316 373316 335368
rect 399024 335316 399076 335368
rect 400864 335316 400916 335368
rect 427360 335316 427412 335368
rect 428464 335316 428516 335368
rect 455328 335316 455380 335368
rect 456064 335316 456116 335368
rect 483204 335316 483256 335368
rect 485044 335316 485096 335368
rect 511356 335316 511408 335368
rect 512644 335316 512696 335368
rect 539324 335316 539376 335368
rect 540244 335316 540296 335368
rect 567200 335316 567252 335368
rect 37924 333208 37976 333260
rect 545764 333208 545816 333260
rect 35624 332528 35676 332580
rect 36820 332528 36872 332580
rect 209688 331236 209740 331288
rect 262220 331236 262272 331288
rect 266268 331236 266320 331288
rect 317420 331236 317472 331288
rect 405648 331236 405700 331288
rect 458180 331236 458232 331288
rect 462228 331236 462280 331288
rect 513380 331236 513432 331288
rect 483664 315936 483716 315988
rect 491668 315936 491720 315988
rect 428648 315256 428700 315308
rect 435732 315256 435784 315308
rect 512736 315256 512788 315308
rect 519636 315256 519688 315308
rect 232688 315120 232740 315172
rect 239772 315120 239824 315172
rect 63592 314644 63644 314696
rect 64328 314644 64380 314696
rect 287704 314644 287756 314696
rect 295708 314644 295760 314696
rect 316776 314644 316828 314696
rect 323676 314644 323728 314696
rect 13728 314576 13780 314628
rect 66260 314576 66312 314628
rect 70308 314576 70360 314628
rect 121460 314576 121512 314628
rect 126888 314576 126940 314628
rect 178040 314576 178092 314628
rect 182088 314576 182140 314628
rect 233240 314576 233292 314628
rect 238668 314576 238720 314628
rect 289820 314576 289872 314628
rect 293868 314576 293920 314628
rect 345020 314576 345072 314628
rect 350448 314576 350500 314628
rect 401600 314576 401652 314628
rect 427728 314576 427780 314628
rect 428556 314576 428608 314628
rect 434628 314576 434680 314628
rect 485780 314576 485832 314628
rect 489828 314576 489880 314628
rect 542360 314576 542412 314628
rect 35624 314508 35676 314560
rect 37004 314508 37056 314560
rect 42708 314508 42760 314560
rect 93860 314508 93912 314560
rect 97908 314508 97960 314560
rect 149060 314508 149112 314560
rect 154488 314508 154540 314560
rect 205640 314508 205692 314560
rect 259736 314508 259788 314560
rect 260196 314508 260248 314560
rect 322848 314508 322900 314560
rect 374000 314508 374052 314560
rect 378048 314508 378100 314560
rect 429200 314508 429252 314560
rect 455696 314508 455748 314560
rect 456156 314508 456208 314560
rect 518808 314508 518860 314560
rect 569960 314508 570012 314560
rect 343548 314440 343600 314492
rect 345664 314440 345716 314492
rect 25688 311788 25740 311840
rect 36728 311788 36780 311840
rect 42892 311788 42944 311840
rect 15200 311720 15252 311772
rect 43996 311720 44048 311772
rect 72056 311788 72108 311840
rect 99472 311788 99524 311840
rect 71872 311720 71924 311772
rect 100024 311720 100076 311772
rect 127072 311788 127124 311840
rect 127992 311720 128044 311772
rect 183652 311788 183704 311840
rect 156052 311720 156104 311772
rect 165988 311720 166040 311772
rect 177304 311720 177356 311772
rect 178684 311720 178736 311772
rect 184020 311720 184072 311772
rect 374644 311788 374696 311840
rect 379704 311788 379756 311840
rect 539324 311788 539376 311840
rect 543004 311788 543056 311840
rect 211712 311720 211764 311772
rect 222016 311720 222068 311772
rect 232596 311720 232648 311772
rect 249708 311720 249760 311772
rect 260104 311720 260156 311772
rect 261484 311720 261536 311772
rect 567200 311720 567252 311772
rect 53656 311652 53708 311704
rect 69664 311652 69716 311704
rect 81992 311652 82044 311704
rect 94504 311652 94556 311704
rect 109684 311652 109736 311704
rect 120724 311652 120776 311704
rect 137652 311652 137704 311704
rect 148416 311652 148468 311704
rect 193680 311652 193732 311704
rect 204904 311652 204956 311704
rect 238852 311652 238904 311704
rect 268016 311652 268068 311704
rect 277676 311652 277728 311704
rect 289084 311652 289136 311704
rect 306012 311652 306064 311704
rect 316684 311652 316736 311704
rect 323032 311652 323084 311704
rect 352012 311652 352064 311704
rect 361672 311652 361724 311704
rect 373264 311652 373316 311704
rect 379612 311652 379664 311704
rect 408040 311652 408092 311704
rect 417700 311652 417752 311704
rect 428464 311652 428516 311704
rect 434812 311652 434864 311704
rect 463700 311652 463752 311704
rect 474004 311652 474056 311704
rect 485044 311652 485096 311704
rect 501696 311652 501748 311704
rect 512644 311652 512696 311704
rect 518992 311652 519044 311704
rect 547880 311652 547932 311704
rect 333704 311584 333756 311636
rect 344284 311584 344336 311636
rect 390008 311584 390060 311636
rect 400864 311584 400916 311636
rect 445668 311584 445720 311636
rect 456064 311584 456116 311636
rect 529664 311584 529716 311636
rect 540244 311584 540296 311636
rect 36912 311516 36964 311568
rect 557540 311516 557592 311568
rect 16028 308388 16080 308440
rect 547880 308388 547932 308440
rect 25688 308048 25740 308100
rect 261484 308048 261536 308100
rect 148324 307980 148376 308032
rect 165620 307980 165672 308032
rect 175464 307980 175516 308032
rect 193680 307980 193732 308032
rect 203524 307980 203576 308032
rect 221372 307980 221424 308032
rect 296352 307980 296404 308032
rect 316776 307980 316828 308032
rect 408040 307980 408092 308032
rect 428648 307980 428700 308032
rect 492036 307980 492088 308032
rect 512736 307980 512788 308032
rect 37004 307912 37056 307964
rect 53656 307912 53708 307964
rect 64328 307912 64380 307964
rect 81440 307912 81492 307964
rect 91468 307912 91520 307964
rect 109684 307912 109736 307964
rect 119436 307912 119488 307964
rect 137652 307912 137704 307964
rect 156328 307912 156380 307964
rect 178684 307912 178736 307964
rect 232596 307912 232648 307964
rect 249708 307912 249760 307964
rect 260196 307912 260248 307964
rect 277676 307912 277728 307964
rect 287520 307912 287572 307964
rect 305368 307912 305420 307964
rect 345664 307912 345716 307964
rect 361672 307912 361724 307964
rect 371516 307912 371568 307964
rect 389364 307912 389416 307964
rect 399484 307912 399536 307964
rect 417700 307912 417752 307964
rect 456064 307912 456116 307964
rect 473544 307912 473596 307964
rect 483480 307912 483532 307964
rect 501696 307912 501748 307964
rect 36912 307844 36964 307896
rect 63316 307844 63368 307896
rect 66904 307844 66956 307896
rect 91100 307844 91152 307896
rect 94504 307844 94556 307896
rect 119344 307844 119396 307896
rect 120724 307844 120776 307896
rect 147312 307844 147364 307896
rect 148416 307844 148468 307896
rect 175280 307844 175332 307896
rect 177304 307844 177356 307896
rect 203340 307844 203392 307896
rect 204904 307844 204956 307896
rect 231032 307844 231084 307896
rect 232504 307844 232556 307896
rect 259368 307844 259420 307896
rect 268016 307844 268068 307896
rect 287704 307844 287756 307896
rect 315488 307844 315540 307896
rect 333704 307844 333756 307896
rect 352012 307844 352064 307896
rect 374644 307844 374696 307896
rect 428556 307844 428608 307896
rect 445668 307844 445720 307896
rect 464344 307844 464396 307896
rect 483664 307844 483716 307896
rect 511448 307844 511500 307896
rect 529664 307844 529716 307896
rect 543004 307844 543056 307896
rect 557540 307844 557592 307896
rect 212264 307776 212316 307828
rect 232688 307776 232740 307828
rect 260104 307776 260156 307828
rect 287336 307776 287388 307828
rect 289084 307776 289136 307828
rect 315028 307776 315080 307828
rect 316684 307776 316736 307828
rect 343364 307776 343416 307828
rect 344284 307776 344336 307828
rect 371332 307776 371384 307828
rect 373264 307776 373316 307828
rect 399024 307776 399076 307828
rect 400864 307776 400916 307828
rect 427360 307776 427412 307828
rect 428464 307776 428516 307828
rect 455328 307776 455380 307828
rect 456156 307776 456208 307828
rect 483204 307776 483256 307828
rect 485044 307776 485096 307828
rect 511356 307776 511408 307828
rect 512644 307776 512696 307828
rect 539324 307776 539376 307828
rect 540244 307776 540296 307828
rect 567200 307776 567252 307828
rect 37924 305600 37976 305652
rect 545764 305600 545816 305652
rect 3056 304988 3108 305040
rect 10324 304988 10376 305040
rect 35624 304988 35676 305040
rect 36728 304988 36780 305040
rect 63592 291864 63644 291916
rect 64328 291864 64380 291916
rect 259736 291864 259788 291916
rect 260196 291864 260248 291916
rect 287704 288328 287756 288380
rect 295708 288328 295760 288380
rect 316776 288328 316828 288380
rect 323676 288328 323728 288380
rect 232688 287920 232740 287972
rect 239772 287920 239824 287972
rect 428648 287648 428700 287700
rect 435732 287648 435784 287700
rect 512736 287512 512788 287564
rect 519636 287512 519688 287564
rect 483664 287376 483716 287428
rect 491668 287376 491720 287428
rect 13728 286968 13780 287020
rect 66260 286968 66312 287020
rect 70308 286968 70360 287020
rect 121460 286968 121512 287020
rect 126888 286968 126940 287020
rect 178040 286968 178092 287020
rect 209688 286968 209740 287020
rect 262220 286968 262272 287020
rect 266268 286968 266320 287020
rect 317420 286968 317472 287020
rect 322848 286968 322900 287020
rect 374000 286968 374052 287020
rect 405648 286968 405700 287020
rect 458180 286968 458232 287020
rect 489828 286968 489880 287020
rect 542360 286968 542412 287020
rect 35624 286900 35676 286952
rect 37004 286900 37056 286952
rect 42708 286900 42760 286952
rect 93860 286900 93912 286952
rect 97908 286900 97960 286952
rect 149060 286900 149112 286952
rect 154488 286900 154540 286952
rect 205640 286900 205692 286952
rect 238668 286900 238720 286952
rect 289820 286900 289872 286952
rect 293868 286900 293920 286952
rect 182088 286832 182140 286884
rect 233240 286832 233292 286884
rect 343548 286900 343600 286952
rect 345664 286900 345716 286952
rect 350448 286900 350500 286952
rect 401600 286900 401652 286952
rect 434628 286900 434680 286952
rect 485780 286900 485832 286952
rect 518808 286900 518860 286952
rect 569960 286900 570012 286952
rect 345020 286832 345072 286884
rect 378048 286832 378100 286884
rect 429200 286832 429252 286884
rect 462228 286832 462280 286884
rect 513380 286832 513432 286884
rect 231676 286764 231728 286816
rect 232596 286764 232648 286816
rect 427728 286764 427780 286816
rect 428556 286764 428608 286816
rect 539508 286764 539560 286816
rect 543004 286764 543056 286816
rect 25688 284248 25740 284300
rect 36912 284248 36964 284300
rect 178684 284248 178736 284300
rect 184020 284248 184072 284300
rect 374644 284248 374696 284300
rect 379704 284248 379756 284300
rect 15200 284180 15252 284232
rect 43996 284180 44048 284232
rect 71044 284180 71096 284232
rect 567200 284180 567252 284232
rect 53656 284112 53708 284164
rect 66904 284112 66956 284164
rect 71872 284112 71924 284164
rect 100024 284112 100076 284164
rect 42892 284044 42944 284096
rect 72056 284044 72108 284096
rect 81992 284044 82044 284096
rect 94504 284044 94556 284096
rect 99472 284044 99524 284096
rect 127992 284112 128044 284164
rect 109684 284044 109736 284096
rect 120724 284044 120776 284096
rect 127072 284044 127124 284096
rect 156052 284112 156104 284164
rect 165988 284112 166040 284164
rect 177304 284112 177356 284164
rect 183652 284112 183704 284164
rect 211712 284112 211764 284164
rect 222016 284112 222068 284164
rect 232504 284112 232556 284164
rect 238852 284112 238904 284164
rect 268016 284112 268068 284164
rect 277676 284112 277728 284164
rect 289084 284112 289136 284164
rect 306012 284112 306064 284164
rect 316684 284112 316736 284164
rect 323032 284112 323084 284164
rect 352012 284112 352064 284164
rect 361672 284112 361724 284164
rect 373264 284112 373316 284164
rect 379612 284112 379664 284164
rect 408040 284112 408092 284164
rect 417700 284112 417752 284164
rect 428464 284112 428516 284164
rect 434812 284112 434864 284164
rect 463700 284112 463752 284164
rect 474004 284112 474056 284164
rect 485044 284112 485096 284164
rect 501696 284112 501748 284164
rect 512644 284112 512696 284164
rect 518992 284112 519044 284164
rect 547880 284112 547932 284164
rect 137652 284044 137704 284096
rect 148416 284044 148468 284096
rect 193680 284044 193732 284096
rect 204904 284044 204956 284096
rect 249708 284044 249760 284096
rect 260104 284044 260156 284096
rect 333704 284044 333756 284096
rect 344284 284044 344336 284096
rect 390008 284044 390060 284096
rect 400864 284044 400916 284096
rect 445668 284044 445720 284096
rect 456156 284044 456208 284096
rect 529664 284044 529716 284096
rect 540244 284044 540296 284096
rect 36820 283976 36872 284028
rect 557540 283976 557592 284028
rect 16028 280780 16080 280832
rect 547880 280780 547932 280832
rect 25688 280372 25740 280424
rect 71044 280372 71096 280424
rect 212356 280372 212408 280424
rect 232688 280372 232740 280424
rect 296352 280372 296404 280424
rect 316776 280372 316828 280424
rect 408040 280372 408092 280424
rect 428648 280372 428700 280424
rect 492036 280372 492088 280424
rect 512736 280372 512788 280424
rect 37004 280304 37056 280356
rect 53656 280304 53708 280356
rect 148416 280304 148468 280356
rect 165712 280304 165764 280356
rect 175464 280304 175516 280356
rect 193680 280304 193732 280356
rect 203524 280304 203576 280356
rect 221372 280304 221424 280356
rect 260104 280304 260156 280356
rect 277676 280304 277728 280356
rect 287520 280304 287572 280356
rect 305368 280304 305420 280356
rect 345664 280304 345716 280356
rect 361672 280304 361724 280356
rect 371516 280304 371568 280356
rect 389364 280304 389416 280356
rect 399484 280304 399536 280356
rect 417700 280304 417752 280356
rect 456156 280304 456208 280356
rect 473360 280304 473412 280356
rect 483480 280304 483532 280356
rect 501696 280304 501748 280356
rect 36912 280236 36964 280288
rect 63316 280236 63368 280288
rect 64328 280236 64380 280288
rect 81440 280236 81492 280288
rect 91468 280236 91520 280288
rect 109684 280236 109736 280288
rect 119436 280236 119488 280288
rect 137652 280236 137704 280288
rect 156328 280236 156380 280288
rect 178684 280236 178736 280288
rect 232504 280236 232556 280288
rect 249708 280236 249760 280288
rect 268016 280236 268068 280288
rect 287704 280236 287756 280288
rect 315488 280236 315540 280288
rect 333704 280236 333756 280288
rect 352012 280236 352064 280288
rect 374644 280236 374696 280288
rect 428464 280236 428516 280288
rect 445668 280236 445720 280288
rect 464344 280236 464396 280288
rect 483664 280236 483716 280288
rect 511448 280236 511500 280288
rect 529664 280236 529716 280288
rect 543004 280236 543056 280288
rect 557540 280236 557592 280288
rect 69664 280168 69716 280220
rect 91100 280168 91152 280220
rect 94504 280168 94556 280220
rect 119344 280168 119396 280220
rect 120724 280168 120776 280220
rect 147312 280168 147364 280220
rect 148324 280168 148376 280220
rect 175372 280168 175424 280220
rect 177304 280168 177356 280220
rect 203340 280168 203392 280220
rect 204904 280168 204956 280220
rect 231032 280168 231084 280220
rect 232596 280168 232648 280220
rect 259368 280168 259420 280220
rect 260196 280168 260248 280220
rect 287336 280168 287388 280220
rect 289084 280168 289136 280220
rect 315028 280168 315080 280220
rect 316684 280168 316736 280220
rect 343364 280168 343416 280220
rect 344284 280168 344336 280220
rect 371332 280168 371384 280220
rect 373264 280168 373316 280220
rect 399024 280168 399076 280220
rect 400864 280168 400916 280220
rect 427360 280168 427412 280220
rect 428556 280168 428608 280220
rect 455328 280168 455380 280220
rect 456064 280168 456116 280220
rect 483020 280168 483072 280220
rect 485044 280168 485096 280220
rect 511356 280168 511408 280220
rect 512644 280168 512696 280220
rect 539324 280168 539376 280220
rect 540244 280168 540296 280220
rect 567200 280168 567252 280220
rect 37924 279420 37976 279472
rect 545764 279420 545816 279472
rect 182088 277516 182140 277568
rect 233240 277516 233292 277568
rect 378048 277516 378100 277568
rect 429200 277516 429252 277568
rect 462228 277516 462280 277568
rect 513380 277516 513432 277568
rect 35624 277448 35676 277500
rect 36820 277448 36872 277500
rect 42708 277448 42760 277500
rect 93860 277448 93912 277500
rect 97908 277448 97960 277500
rect 149060 277448 149112 277500
rect 154488 277448 154540 277500
rect 205640 277448 205692 277500
rect 238668 277448 238720 277500
rect 289820 277448 289872 277500
rect 293868 277448 293920 277500
rect 345020 277448 345072 277500
rect 350448 277448 350500 277500
rect 401600 277448 401652 277500
rect 434628 277448 434680 277500
rect 485780 277448 485832 277500
rect 518808 277448 518860 277500
rect 569960 277448 570012 277500
rect 13728 277380 13780 277432
rect 66260 277380 66312 277432
rect 70308 277380 70360 277432
rect 121460 277380 121512 277432
rect 126888 277380 126940 277432
rect 178040 277380 178092 277432
rect 209688 277380 209740 277432
rect 262220 277380 262272 277432
rect 266268 277380 266320 277432
rect 317420 277380 317472 277432
rect 322848 277380 322900 277432
rect 374000 277380 374052 277432
rect 405648 277380 405700 277432
rect 458180 277380 458232 277432
rect 489828 277380 489880 277432
rect 542360 277380 542412 277432
rect 63592 263440 63644 263492
rect 64328 263440 64380 263492
rect 455696 263440 455748 263492
rect 456156 263440 456208 263492
rect 232688 262148 232740 262200
rect 239772 262148 239824 262200
rect 483664 262148 483716 262200
rect 491668 262148 491720 262200
rect 512736 262148 512788 262200
rect 519636 262148 519688 262200
rect 428648 261468 428700 261520
rect 435732 261468 435784 261520
rect 316776 261400 316828 261452
rect 323676 261400 323728 261452
rect 287704 261264 287756 261316
rect 295708 261264 295760 261316
rect 147680 259428 147732 259480
rect 148416 259428 148468 259480
rect 35624 259360 35676 259412
rect 37004 259360 37056 259412
rect 343640 259360 343692 259412
rect 345664 259360 345716 259412
rect 42892 256640 42944 256692
rect 15200 256572 15252 256624
rect 43996 256572 44048 256624
rect 71964 256640 72016 256692
rect 99472 256640 99524 256692
rect 71872 256572 71924 256624
rect 100024 256572 100076 256624
rect 127072 256640 127124 256692
rect 127992 256572 128044 256624
rect 183652 256640 183704 256692
rect 155960 256572 156012 256624
rect 165988 256572 166040 256624
rect 177304 256572 177356 256624
rect 178684 256572 178736 256624
rect 184020 256572 184072 256624
rect 374644 256640 374696 256692
rect 379704 256640 379756 256692
rect 539324 256640 539376 256692
rect 543004 256640 543056 256692
rect 211712 256572 211764 256624
rect 221924 256572 221976 256624
rect 232596 256572 232648 256624
rect 249708 256572 249760 256624
rect 260196 256572 260248 256624
rect 261484 256572 261536 256624
rect 567200 256572 567252 256624
rect 25688 256504 25740 256556
rect 36912 256504 36964 256556
rect 53656 256504 53708 256556
rect 69664 256504 69716 256556
rect 81992 256504 82044 256556
rect 94504 256504 94556 256556
rect 109684 256504 109736 256556
rect 120724 256504 120776 256556
rect 137652 256504 137704 256556
rect 148324 256504 148376 256556
rect 193680 256504 193732 256556
rect 204904 256504 204956 256556
rect 238852 256504 238904 256556
rect 268016 256504 268068 256556
rect 277676 256504 277728 256556
rect 289084 256504 289136 256556
rect 306012 256504 306064 256556
rect 316684 256504 316736 256556
rect 323032 256504 323084 256556
rect 352012 256504 352064 256556
rect 361672 256504 361724 256556
rect 373264 256504 373316 256556
rect 379612 256504 379664 256556
rect 408040 256504 408092 256556
rect 417700 256504 417752 256556
rect 428556 256504 428608 256556
rect 434812 256504 434864 256556
rect 463792 256504 463844 256556
rect 474004 256504 474056 256556
rect 485044 256504 485096 256556
rect 501696 256504 501748 256556
rect 512644 256504 512696 256556
rect 518992 256504 519044 256556
rect 547880 256504 547932 256556
rect 333704 256436 333756 256488
rect 344284 256436 344336 256488
rect 390008 256436 390060 256488
rect 400864 256436 400916 256488
rect 445668 256436 445720 256488
rect 456064 256436 456116 256488
rect 529664 256436 529716 256488
rect 540244 256436 540296 256488
rect 36728 256368 36780 256420
rect 557540 256368 557592 256420
rect 16028 254532 16080 254584
rect 547880 254532 547932 254584
rect 25688 254124 25740 254176
rect 69664 254124 69716 254176
rect 212356 254124 212408 254176
rect 232688 254124 232740 254176
rect 296352 254124 296404 254176
rect 316776 254124 316828 254176
rect 492036 254124 492088 254176
rect 512736 254124 512788 254176
rect 3332 254056 3384 254108
rect 7656 254056 7708 254108
rect 37004 254056 37056 254108
rect 53656 254056 53708 254108
rect 64328 254056 64380 254108
rect 81440 254056 81492 254108
rect 148416 254056 148468 254108
rect 165712 254056 165764 254108
rect 175464 254056 175516 254108
rect 193680 254056 193732 254108
rect 203524 254056 203576 254108
rect 221372 254056 221424 254108
rect 260196 254056 260248 254108
rect 277676 254056 277728 254108
rect 287520 254056 287572 254108
rect 305368 254056 305420 254108
rect 345664 254056 345716 254108
rect 361672 254056 361724 254108
rect 371516 254056 371568 254108
rect 389364 254056 389416 254108
rect 399484 254056 399536 254108
rect 417700 254056 417752 254108
rect 428556 254056 428608 254108
rect 445668 254056 445720 254108
rect 456064 254056 456116 254108
rect 473360 254056 473412 254108
rect 483480 254056 483532 254108
rect 501696 254056 501748 254108
rect 36912 253988 36964 254040
rect 63316 253988 63368 254040
rect 66904 253988 66956 254040
rect 91100 253988 91152 254040
rect 91468 253988 91520 254040
rect 109684 253988 109736 254040
rect 119436 253988 119488 254040
rect 137652 253988 137704 254040
rect 156328 253988 156380 254040
rect 178684 253988 178736 254040
rect 232596 253988 232648 254040
rect 249708 253988 249760 254040
rect 268016 253988 268068 254040
rect 287704 253988 287756 254040
rect 315488 253988 315540 254040
rect 333704 253988 333756 254040
rect 352012 253988 352064 254040
rect 374644 253988 374696 254040
rect 408040 253988 408092 254040
rect 428648 253988 428700 254040
rect 464344 253988 464396 254040
rect 483664 253988 483716 254040
rect 511448 253988 511500 254040
rect 529664 253988 529716 254040
rect 543004 253988 543056 254040
rect 557540 253988 557592 254040
rect 94504 253920 94556 253972
rect 119344 253920 119396 253972
rect 120724 253920 120776 253972
rect 147312 253920 147364 253972
rect 148324 253920 148376 253972
rect 175372 253920 175424 253972
rect 177304 253920 177356 253972
rect 203340 253920 203392 253972
rect 204904 253920 204956 253972
rect 231032 253920 231084 253972
rect 232504 253920 232556 253972
rect 259368 253920 259420 253972
rect 260104 253920 260156 253972
rect 287336 253920 287388 253972
rect 289084 253920 289136 253972
rect 315028 253920 315080 253972
rect 316684 253920 316736 253972
rect 343364 253920 343416 253972
rect 344284 253920 344336 253972
rect 371332 253920 371384 253972
rect 373264 253920 373316 253972
rect 399024 253920 399076 253972
rect 400864 253920 400916 253972
rect 427360 253920 427412 253972
rect 428464 253920 428516 253972
rect 455328 253920 455380 253972
rect 456156 253920 456208 253972
rect 483020 253920 483072 253972
rect 485044 253920 485096 253972
rect 511356 253920 511408 253972
rect 512644 253920 512696 253972
rect 539324 253920 539376 253972
rect 540244 253920 540296 253972
rect 567200 253920 567252 253972
rect 37924 251812 37976 251864
rect 545764 251812 545816 251864
rect 182088 251268 182140 251320
rect 233240 251268 233292 251320
rect 378048 251268 378100 251320
rect 429200 251268 429252 251320
rect 35624 251200 35676 251252
rect 36728 251200 36780 251252
rect 42708 251200 42760 251252
rect 93860 251200 93912 251252
rect 97908 251200 97960 251252
rect 149060 251200 149112 251252
rect 154488 251200 154540 251252
rect 205640 251200 205692 251252
rect 238668 251200 238720 251252
rect 289820 251200 289872 251252
rect 293868 251200 293920 251252
rect 345020 251200 345072 251252
rect 350448 251200 350500 251252
rect 401600 251200 401652 251252
rect 434628 251200 434680 251252
rect 485780 251200 485832 251252
rect 489828 251200 489880 251252
rect 542360 251200 542412 251252
rect 3056 240184 3108 240236
rect 6276 240184 6328 240236
rect 63592 235356 63644 235408
rect 64328 235356 64380 235408
rect 147680 235356 147732 235408
rect 148416 235356 148468 235408
rect 259736 235356 259788 235408
rect 260196 235356 260248 235408
rect 512736 234200 512788 234252
rect 519636 234200 519688 234252
rect 428648 233860 428700 233912
rect 435732 233860 435784 233912
rect 232688 233520 232740 233572
rect 239772 233520 239824 233572
rect 287704 233520 287756 233572
rect 295708 233520 295760 233572
rect 316776 233384 316828 233436
rect 323676 233384 323728 233436
rect 483664 233384 483716 233436
rect 491668 233384 491720 233436
rect 13728 233180 13780 233232
rect 66260 233180 66312 233232
rect 70308 233180 70360 233232
rect 121460 233180 121512 233232
rect 126888 233180 126940 233232
rect 178040 233180 178092 233232
rect 209688 233180 209740 233232
rect 262220 233180 262272 233232
rect 266268 233180 266320 233232
rect 317420 233180 317472 233232
rect 322848 233180 322900 233232
rect 374000 233180 374052 233232
rect 405648 233180 405700 233232
rect 458180 233180 458232 233232
rect 462228 233180 462280 233232
rect 513380 233180 513432 233232
rect 518808 233180 518860 233232
rect 569960 233180 570012 233232
rect 231676 233112 231728 233164
rect 232596 233112 232648 233164
rect 427728 233112 427780 233164
rect 428556 233112 428608 233164
rect 539508 233112 539560 233164
rect 543004 233112 543056 233164
rect 35624 232704 35676 232756
rect 37004 232704 37056 232756
rect 343640 232704 343692 232756
rect 345664 232704 345716 232756
rect 178684 230392 178736 230444
rect 184020 230392 184072 230444
rect 374644 230392 374696 230444
rect 379704 230392 379756 230444
rect 15200 230324 15252 230376
rect 43996 230324 44048 230376
rect 71044 230324 71096 230376
rect 567200 230324 567252 230376
rect 25688 230256 25740 230308
rect 36912 230256 36964 230308
rect 53656 230256 53708 230308
rect 66904 230256 66956 230308
rect 71872 230256 71924 230308
rect 100024 230256 100076 230308
rect 42892 230188 42944 230240
rect 72056 230188 72108 230240
rect 81992 230188 82044 230240
rect 94504 230188 94556 230240
rect 99472 230188 99524 230240
rect 127992 230256 128044 230308
rect 109684 230188 109736 230240
rect 120724 230188 120776 230240
rect 127072 230188 127124 230240
rect 156052 230256 156104 230308
rect 165988 230256 166040 230308
rect 177304 230256 177356 230308
rect 183652 230256 183704 230308
rect 211712 230256 211764 230308
rect 222016 230256 222068 230308
rect 232504 230256 232556 230308
rect 238852 230256 238904 230308
rect 268016 230256 268068 230308
rect 277676 230256 277728 230308
rect 289084 230256 289136 230308
rect 306012 230256 306064 230308
rect 316684 230256 316736 230308
rect 323032 230256 323084 230308
rect 352012 230256 352064 230308
rect 361672 230256 361724 230308
rect 373264 230256 373316 230308
rect 379612 230256 379664 230308
rect 408040 230256 408092 230308
rect 417700 230256 417752 230308
rect 428464 230256 428516 230308
rect 434812 230256 434864 230308
rect 463700 230256 463752 230308
rect 474004 230256 474056 230308
rect 485044 230256 485096 230308
rect 501696 230256 501748 230308
rect 512644 230256 512696 230308
rect 518992 230256 519044 230308
rect 547880 230256 547932 230308
rect 137652 230188 137704 230240
rect 148324 230188 148376 230240
rect 193680 230188 193732 230240
rect 204904 230188 204956 230240
rect 249708 230188 249760 230240
rect 260104 230188 260156 230240
rect 333704 230188 333756 230240
rect 344284 230188 344336 230240
rect 390008 230188 390060 230240
rect 400864 230188 400916 230240
rect 445668 230188 445720 230240
rect 456156 230188 456208 230240
rect 529664 230188 529716 230240
rect 540244 230188 540296 230240
rect 36820 230120 36872 230172
rect 557540 230120 557592 230172
rect 15292 226992 15344 227044
rect 547880 226992 547932 227044
rect 25688 226584 25740 226636
rect 261484 226584 261536 226636
rect 148324 226516 148376 226568
rect 165712 226516 165764 226568
rect 175464 226516 175516 226568
rect 193680 226516 193732 226568
rect 203524 226516 203576 226568
rect 221372 226516 221424 226568
rect 296352 226516 296404 226568
rect 316776 226516 316828 226568
rect 408040 226516 408092 226568
rect 428648 226516 428700 226568
rect 492036 226516 492088 226568
rect 512736 226516 512788 226568
rect 37004 226448 37056 226500
rect 53656 226448 53708 226500
rect 64328 226448 64380 226500
rect 81440 226448 81492 226500
rect 91468 226448 91520 226500
rect 109684 226448 109736 226500
rect 119436 226448 119488 226500
rect 137652 226448 137704 226500
rect 156328 226448 156380 226500
rect 178684 226448 178736 226500
rect 232504 226448 232556 226500
rect 249708 226448 249760 226500
rect 260196 226448 260248 226500
rect 277676 226448 277728 226500
rect 287520 226448 287572 226500
rect 305368 226448 305420 226500
rect 345664 226448 345716 226500
rect 361672 226448 361724 226500
rect 371516 226448 371568 226500
rect 389364 226448 389416 226500
rect 399484 226448 399536 226500
rect 417700 226448 417752 226500
rect 456156 226448 456208 226500
rect 473360 226448 473412 226500
rect 483480 226448 483532 226500
rect 501696 226448 501748 226500
rect 36912 226380 36964 226432
rect 63316 226380 63368 226432
rect 66904 226380 66956 226432
rect 91100 226380 91152 226432
rect 94504 226380 94556 226432
rect 119344 226380 119396 226432
rect 120724 226380 120776 226432
rect 147312 226380 147364 226432
rect 148416 226380 148468 226432
rect 175372 226380 175424 226432
rect 177304 226380 177356 226432
rect 203340 226380 203392 226432
rect 204904 226380 204956 226432
rect 231032 226380 231084 226432
rect 232596 226380 232648 226432
rect 259368 226380 259420 226432
rect 268016 226380 268068 226432
rect 287704 226380 287756 226432
rect 315488 226380 315540 226432
rect 333704 226380 333756 226432
rect 352012 226380 352064 226432
rect 374644 226380 374696 226432
rect 428556 226380 428608 226432
rect 445668 226380 445720 226432
rect 464344 226380 464396 226432
rect 483664 226380 483716 226432
rect 511448 226380 511500 226432
rect 529664 226380 529716 226432
rect 543004 226380 543056 226432
rect 557540 226380 557592 226432
rect 212356 226312 212408 226364
rect 232688 226312 232740 226364
rect 260104 226312 260156 226364
rect 287336 226312 287388 226364
rect 289084 226312 289136 226364
rect 315028 226312 315080 226364
rect 316684 226312 316736 226364
rect 343364 226312 343416 226364
rect 344284 226312 344336 226364
rect 371332 226312 371384 226364
rect 373264 226312 373316 226364
rect 399024 226312 399076 226364
rect 400864 226312 400916 226364
rect 427360 226312 427412 226364
rect 428464 226312 428516 226364
rect 455328 226312 455380 226364
rect 456064 226312 456116 226364
rect 483020 226312 483072 226364
rect 485044 226312 485096 226364
rect 511356 226312 511408 226364
rect 512644 226312 512696 226364
rect 539324 226312 539376 226364
rect 540244 226312 540296 226364
rect 567200 226312 567252 226364
rect 37924 225564 37976 225616
rect 545764 225564 545816 225616
rect 35624 223592 35676 223644
rect 36820 223592 36872 223644
rect 232688 207748 232740 207800
rect 239772 207748 239824 207800
rect 428648 207612 428700 207664
rect 435732 207612 435784 207664
rect 483664 207408 483716 207460
rect 491668 207408 491720 207460
rect 63592 207340 63644 207392
rect 64328 207340 64380 207392
rect 259736 207340 259788 207392
rect 260196 207340 260248 207392
rect 316776 207340 316828 207392
rect 323676 207340 323728 207392
rect 455696 207340 455748 207392
rect 456156 207340 456208 207392
rect 512736 207272 512788 207324
rect 519636 207272 519688 207324
rect 287704 207136 287756 207188
rect 295708 207136 295760 207188
rect 13728 205572 13780 205624
rect 66260 205572 66312 205624
rect 70308 205572 70360 205624
rect 121460 205572 121512 205624
rect 126888 205572 126940 205624
rect 178040 205572 178092 205624
rect 209688 205572 209740 205624
rect 262220 205572 262272 205624
rect 266268 205572 266320 205624
rect 317420 205572 317472 205624
rect 322848 205572 322900 205624
rect 374000 205572 374052 205624
rect 405648 205572 405700 205624
rect 458180 205572 458232 205624
rect 489828 205572 489880 205624
rect 542360 205572 542412 205624
rect 35624 205504 35676 205556
rect 37004 205504 37056 205556
rect 42708 205504 42760 205556
rect 93860 205504 93912 205556
rect 97908 205504 97960 205556
rect 149060 205504 149112 205556
rect 154488 205504 154540 205556
rect 205640 205504 205692 205556
rect 238668 205504 238720 205556
rect 289820 205504 289872 205556
rect 293868 205504 293920 205556
rect 345020 205504 345072 205556
rect 350448 205504 350500 205556
rect 401600 205504 401652 205556
rect 427728 205504 427780 205556
rect 428556 205504 428608 205556
rect 434628 205504 434680 205556
rect 485780 205504 485832 205556
rect 518808 205504 518860 205556
rect 569960 205504 570012 205556
rect 182088 205436 182140 205488
rect 233240 205436 233292 205488
rect 343640 205436 343692 205488
rect 345664 205436 345716 205488
rect 378048 205436 378100 205488
rect 429200 205436 429252 205488
rect 462228 205436 462280 205488
rect 513380 205436 513432 205488
rect 539508 205436 539560 205488
rect 543004 205436 543056 205488
rect 178684 202784 178736 202836
rect 184020 202784 184072 202836
rect 374644 202784 374696 202836
rect 379704 202784 379756 202836
rect 15200 202716 15252 202768
rect 43628 202716 43680 202768
rect 69664 202716 69716 202768
rect 567200 202716 567252 202768
rect 25688 202648 25740 202700
rect 36912 202648 36964 202700
rect 53564 202648 53616 202700
rect 66904 202648 66956 202700
rect 71872 202648 71924 202700
rect 100024 202648 100076 202700
rect 42892 202580 42944 202632
rect 72056 202580 72108 202632
rect 81992 202580 82044 202632
rect 94504 202580 94556 202632
rect 99472 202580 99524 202632
rect 127716 202648 127768 202700
rect 109684 202580 109736 202632
rect 120724 202580 120776 202632
rect 127072 202580 127124 202632
rect 156052 202648 156104 202700
rect 165988 202648 166040 202700
rect 177304 202648 177356 202700
rect 183652 202648 183704 202700
rect 211712 202648 211764 202700
rect 222016 202648 222068 202700
rect 232596 202648 232648 202700
rect 238852 202648 238904 202700
rect 268016 202648 268068 202700
rect 277676 202648 277728 202700
rect 289084 202648 289136 202700
rect 306012 202648 306064 202700
rect 316684 202648 316736 202700
rect 323032 202648 323084 202700
rect 352012 202648 352064 202700
rect 361672 202648 361724 202700
rect 373264 202648 373316 202700
rect 379612 202648 379664 202700
rect 408040 202648 408092 202700
rect 417700 202648 417752 202700
rect 428464 202648 428516 202700
rect 434812 202648 434864 202700
rect 463700 202648 463752 202700
rect 474004 202648 474056 202700
rect 485044 202648 485096 202700
rect 501696 202648 501748 202700
rect 512644 202648 512696 202700
rect 518992 202648 519044 202700
rect 547880 202648 547932 202700
rect 137928 202580 137980 202632
rect 148416 202580 148468 202632
rect 193680 202580 193732 202632
rect 204904 202580 204956 202632
rect 249524 202580 249576 202632
rect 260104 202580 260156 202632
rect 333888 202580 333940 202632
rect 344284 202580 344336 202632
rect 390008 202580 390060 202632
rect 400864 202580 400916 202632
rect 445668 202580 445720 202632
rect 456064 202580 456116 202632
rect 529664 202580 529716 202632
rect 540244 202580 540296 202632
rect 36728 202512 36780 202564
rect 557540 202512 557592 202564
rect 16028 200744 16080 200796
rect 547880 200744 547932 200796
rect 25688 200336 25740 200388
rect 71044 200336 71096 200388
rect 212264 200336 212316 200388
rect 232688 200336 232740 200388
rect 296352 200336 296404 200388
rect 316776 200336 316828 200388
rect 408040 200336 408092 200388
rect 428648 200336 428700 200388
rect 492036 200336 492088 200388
rect 512736 200336 512788 200388
rect 36912 200268 36964 200320
rect 53656 200268 53708 200320
rect 148416 200268 148468 200320
rect 165620 200268 165672 200320
rect 175464 200268 175516 200320
rect 193680 200268 193732 200320
rect 203524 200268 203576 200320
rect 221372 200268 221424 200320
rect 260196 200268 260248 200320
rect 277676 200268 277728 200320
rect 287520 200268 287572 200320
rect 305368 200268 305420 200320
rect 345664 200268 345716 200320
rect 361672 200268 361724 200320
rect 371516 200268 371568 200320
rect 389364 200268 389416 200320
rect 399484 200268 399536 200320
rect 417700 200268 417752 200320
rect 456156 200268 456208 200320
rect 473544 200268 473596 200320
rect 483480 200268 483532 200320
rect 501696 200268 501748 200320
rect 37004 200200 37056 200252
rect 63316 200200 63368 200252
rect 64328 200200 64380 200252
rect 81440 200200 81492 200252
rect 91468 200200 91520 200252
rect 109684 200200 109736 200252
rect 119436 200200 119488 200252
rect 137652 200200 137704 200252
rect 156328 200200 156380 200252
rect 178684 200200 178736 200252
rect 232596 200200 232648 200252
rect 249708 200200 249760 200252
rect 268016 200200 268068 200252
rect 287704 200200 287756 200252
rect 315488 200200 315540 200252
rect 333704 200200 333756 200252
rect 352012 200200 352064 200252
rect 374644 200200 374696 200252
rect 428464 200200 428516 200252
rect 445668 200200 445720 200252
rect 464344 200200 464396 200252
rect 483664 200200 483716 200252
rect 511448 200200 511500 200252
rect 529664 200200 529716 200252
rect 543004 200200 543056 200252
rect 557540 200200 557592 200252
rect 69664 200132 69716 200184
rect 91100 200132 91152 200184
rect 94504 200132 94556 200184
rect 119344 200132 119396 200184
rect 120724 200132 120776 200184
rect 147312 200132 147364 200184
rect 148324 200132 148376 200184
rect 175280 200132 175332 200184
rect 177304 200132 177356 200184
rect 203340 200132 203392 200184
rect 204904 200132 204956 200184
rect 231032 200132 231084 200184
rect 232504 200132 232556 200184
rect 259368 200132 259420 200184
rect 260104 200132 260156 200184
rect 287336 200132 287388 200184
rect 289084 200132 289136 200184
rect 315028 200132 315080 200184
rect 316684 200132 316736 200184
rect 343364 200132 343416 200184
rect 344284 200132 344336 200184
rect 371332 200132 371384 200184
rect 373264 200132 373316 200184
rect 399024 200132 399076 200184
rect 400864 200132 400916 200184
rect 427360 200132 427412 200184
rect 428556 200132 428608 200184
rect 455328 200132 455380 200184
rect 456064 200132 456116 200184
rect 483204 200132 483256 200184
rect 485044 200132 485096 200184
rect 511356 200132 511408 200184
rect 512644 200132 512696 200184
rect 539324 200132 539376 200184
rect 540244 200132 540296 200184
rect 567200 200132 567252 200184
rect 37924 197956 37976 198008
rect 545764 197956 545816 198008
rect 35624 197344 35676 197396
rect 36728 197344 36780 197396
rect 2964 187688 3016 187740
rect 13176 187688 13228 187740
rect 63592 185580 63644 185632
rect 64328 185580 64380 185632
rect 147680 185580 147732 185632
rect 148416 185580 148468 185632
rect 259736 185580 259788 185632
rect 260196 185580 260248 185632
rect 455696 185580 455748 185632
rect 456156 185580 456208 185632
rect 428648 180072 428700 180124
rect 435732 180072 435784 180124
rect 232688 179868 232740 179920
rect 239772 179868 239824 179920
rect 512736 179800 512788 179852
rect 519636 179800 519688 179852
rect 483664 179664 483716 179716
rect 491668 179664 491720 179716
rect 287704 179392 287756 179444
rect 295708 179392 295760 179444
rect 316776 179392 316828 179444
rect 323676 179392 323728 179444
rect 13728 179324 13780 179376
rect 66260 179324 66312 179376
rect 70308 179324 70360 179376
rect 121460 179324 121512 179376
rect 126888 179324 126940 179376
rect 178040 179324 178092 179376
rect 209688 179324 209740 179376
rect 262220 179324 262272 179376
rect 266268 179324 266320 179376
rect 317420 179324 317472 179376
rect 322848 179324 322900 179376
rect 374000 179324 374052 179376
rect 405648 179324 405700 179376
rect 458180 179324 458232 179376
rect 489828 179324 489880 179376
rect 542360 179324 542412 179376
rect 35624 179256 35676 179308
rect 36912 179256 36964 179308
rect 42708 179256 42760 179308
rect 93860 179256 93912 179308
rect 97908 179256 97960 179308
rect 149060 179256 149112 179308
rect 154488 179256 154540 179308
rect 205640 179256 205692 179308
rect 231676 179256 231728 179308
rect 232596 179256 232648 179308
rect 238668 179256 238720 179308
rect 289820 179256 289872 179308
rect 293868 179256 293920 179308
rect 182088 179188 182140 179240
rect 233240 179188 233292 179240
rect 343548 179256 343600 179308
rect 345664 179256 345716 179308
rect 350448 179256 350500 179308
rect 401600 179256 401652 179308
rect 434628 179256 434680 179308
rect 485780 179256 485832 179308
rect 518808 179256 518860 179308
rect 569960 179256 570012 179308
rect 345020 179188 345072 179240
rect 378048 179188 378100 179240
rect 429200 179188 429252 179240
rect 462228 179188 462280 179240
rect 513380 179188 513432 179240
rect 42892 176604 42944 176656
rect 15200 176536 15252 176588
rect 43996 176536 44048 176588
rect 72056 176604 72108 176656
rect 99472 176604 99524 176656
rect 71872 176536 71924 176588
rect 100024 176536 100076 176588
rect 127072 176604 127124 176656
rect 127992 176536 128044 176588
rect 183652 176604 183704 176656
rect 156052 176536 156104 176588
rect 165988 176536 166040 176588
rect 177304 176536 177356 176588
rect 178684 176536 178736 176588
rect 184020 176536 184072 176588
rect 374644 176604 374696 176656
rect 379704 176604 379756 176656
rect 539324 176604 539376 176656
rect 543004 176604 543056 176656
rect 211712 176536 211764 176588
rect 222016 176536 222068 176588
rect 232504 176536 232556 176588
rect 249708 176536 249760 176588
rect 260104 176536 260156 176588
rect 261484 176536 261536 176588
rect 567200 176536 567252 176588
rect 25688 176468 25740 176520
rect 37004 176468 37056 176520
rect 53656 176468 53708 176520
rect 69664 176468 69716 176520
rect 81992 176468 82044 176520
rect 94504 176468 94556 176520
rect 109684 176468 109736 176520
rect 120724 176468 120776 176520
rect 137652 176468 137704 176520
rect 148324 176468 148376 176520
rect 193680 176468 193732 176520
rect 204904 176468 204956 176520
rect 238852 176468 238904 176520
rect 268016 176468 268068 176520
rect 277676 176468 277728 176520
rect 289084 176468 289136 176520
rect 306012 176468 306064 176520
rect 316684 176468 316736 176520
rect 323032 176468 323084 176520
rect 352012 176468 352064 176520
rect 361672 176468 361724 176520
rect 373264 176468 373316 176520
rect 379612 176468 379664 176520
rect 408040 176468 408092 176520
rect 417700 176468 417752 176520
rect 428556 176468 428608 176520
rect 434812 176468 434864 176520
rect 463700 176468 463752 176520
rect 474004 176468 474056 176520
rect 485044 176468 485096 176520
rect 501696 176468 501748 176520
rect 512644 176468 512696 176520
rect 518992 176468 519044 176520
rect 547880 176468 547932 176520
rect 333704 176400 333756 176452
rect 344284 176400 344336 176452
rect 390008 176400 390060 176452
rect 400864 176400 400916 176452
rect 445668 176400 445720 176452
rect 456064 176400 456116 176452
rect 529664 176400 529716 176452
rect 540244 176400 540296 176452
rect 36820 176332 36872 176384
rect 557540 176332 557592 176384
rect 16028 173136 16080 173188
rect 547880 173136 547932 173188
rect 212264 172728 212316 172780
rect 232688 172728 232740 172780
rect 296352 172728 296404 172780
rect 316776 172728 316828 172780
rect 408040 172728 408092 172780
rect 428648 172728 428700 172780
rect 492036 172728 492088 172780
rect 512736 172728 512788 172780
rect 25688 172660 25740 172712
rect 39304 172660 39356 172712
rect 148416 172660 148468 172712
rect 165620 172660 165672 172712
rect 175464 172660 175516 172712
rect 193680 172660 193732 172712
rect 203524 172660 203576 172712
rect 221372 172660 221424 172712
rect 260196 172660 260248 172712
rect 277676 172660 277728 172712
rect 287520 172660 287572 172712
rect 305368 172660 305420 172712
rect 345664 172660 345716 172712
rect 361672 172660 361724 172712
rect 371516 172660 371568 172712
rect 389364 172660 389416 172712
rect 399484 172660 399536 172712
rect 417700 172660 417752 172712
rect 456156 172660 456208 172712
rect 473544 172660 473596 172712
rect 483480 172660 483532 172712
rect 501696 172660 501748 172712
rect 37004 172592 37056 172644
rect 53656 172592 53708 172644
rect 64328 172592 64380 172644
rect 81440 172592 81492 172644
rect 91468 172592 91520 172644
rect 109684 172592 109736 172644
rect 119436 172592 119488 172644
rect 137652 172592 137704 172644
rect 156328 172592 156380 172644
rect 178684 172592 178736 172644
rect 232596 172592 232648 172644
rect 249708 172592 249760 172644
rect 268016 172592 268068 172644
rect 287704 172592 287756 172644
rect 315488 172592 315540 172644
rect 333704 172592 333756 172644
rect 352012 172592 352064 172644
rect 374644 172592 374696 172644
rect 428464 172592 428516 172644
rect 445668 172592 445720 172644
rect 464344 172592 464396 172644
rect 483664 172592 483716 172644
rect 511448 172592 511500 172644
rect 529664 172592 529716 172644
rect 543004 172592 543056 172644
rect 557540 172592 557592 172644
rect 36912 172524 36964 172576
rect 63316 172524 63368 172576
rect 66904 172524 66956 172576
rect 91100 172524 91152 172576
rect 94504 172524 94556 172576
rect 119344 172524 119396 172576
rect 120724 172524 120776 172576
rect 147312 172524 147364 172576
rect 148324 172524 148376 172576
rect 175280 172524 175332 172576
rect 177304 172524 177356 172576
rect 203340 172524 203392 172576
rect 204904 172524 204956 172576
rect 231032 172524 231084 172576
rect 232504 172524 232556 172576
rect 259368 172524 259420 172576
rect 260104 172524 260156 172576
rect 287336 172524 287388 172576
rect 289084 172524 289136 172576
rect 315028 172524 315080 172576
rect 316684 172524 316736 172576
rect 343364 172524 343416 172576
rect 344284 172524 344336 172576
rect 371332 172524 371384 172576
rect 373264 172524 373316 172576
rect 399024 172524 399076 172576
rect 400864 172524 400916 172576
rect 427360 172524 427412 172576
rect 428556 172524 428608 172576
rect 455328 172524 455380 172576
rect 456064 172524 456116 172576
rect 483204 172524 483256 172576
rect 485044 172524 485096 172576
rect 511356 172524 511408 172576
rect 512644 172524 512696 172576
rect 539324 172524 539376 172576
rect 540244 172524 540296 172576
rect 567200 172524 567252 172576
rect 37924 170348 37976 170400
rect 545764 170348 545816 170400
rect 35624 169736 35676 169788
rect 36820 169736 36872 169788
rect 63592 156612 63644 156664
rect 64328 156612 64380 156664
rect 147680 156612 147732 156664
rect 148416 156612 148468 156664
rect 259736 156612 259788 156664
rect 260196 156612 260248 156664
rect 455696 156612 455748 156664
rect 456156 156612 456208 156664
rect 287704 153144 287756 153196
rect 295708 153144 295760 153196
rect 316776 153144 316828 153196
rect 323676 153144 323728 153196
rect 232688 152532 232740 152584
rect 239772 152532 239824 152584
rect 428648 152464 428700 152516
rect 435732 152464 435784 152516
rect 483664 152464 483716 152516
rect 491668 152464 491720 152516
rect 512736 152192 512788 152244
rect 519636 152192 519688 152244
rect 13728 151716 13780 151768
rect 66260 151716 66312 151768
rect 70308 151716 70360 151768
rect 121460 151716 121512 151768
rect 126888 151716 126940 151768
rect 178040 151716 178092 151768
rect 209688 151716 209740 151768
rect 262220 151716 262272 151768
rect 266268 151716 266320 151768
rect 317420 151716 317472 151768
rect 322848 151716 322900 151768
rect 374000 151716 374052 151768
rect 405648 151716 405700 151768
rect 458180 151716 458232 151768
rect 489828 151716 489880 151768
rect 542360 151716 542412 151768
rect 35624 151648 35676 151700
rect 37004 151648 37056 151700
rect 42708 151648 42760 151700
rect 93860 151648 93912 151700
rect 97908 151648 97960 151700
rect 149060 151648 149112 151700
rect 154488 151648 154540 151700
rect 205640 151648 205692 151700
rect 231676 151648 231728 151700
rect 232596 151648 232648 151700
rect 238668 151648 238720 151700
rect 289820 151648 289872 151700
rect 293868 151648 293920 151700
rect 182088 151580 182140 151632
rect 233240 151580 233292 151632
rect 343640 151648 343692 151700
rect 345664 151648 345716 151700
rect 350448 151648 350500 151700
rect 401600 151648 401652 151700
rect 434628 151648 434680 151700
rect 485780 151648 485832 151700
rect 518808 151648 518860 151700
rect 569960 151648 570012 151700
rect 345020 151580 345072 151632
rect 378048 151580 378100 151632
rect 429200 151580 429252 151632
rect 462228 151580 462280 151632
rect 513380 151580 513432 151632
rect 539508 151580 539560 151632
rect 543004 151580 543056 151632
rect 178684 148996 178736 149048
rect 184020 148996 184072 149048
rect 374644 148996 374696 149048
rect 379704 148996 379756 149048
rect 15200 148928 15252 148980
rect 43996 148928 44048 148980
rect 71044 148928 71096 148980
rect 567200 148928 567252 148980
rect 25688 148860 25740 148912
rect 36912 148860 36964 148912
rect 53656 148860 53708 148912
rect 66904 148860 66956 148912
rect 71872 148860 71924 148912
rect 100024 148860 100076 148912
rect 42892 148792 42944 148844
rect 72056 148792 72108 148844
rect 81992 148792 82044 148844
rect 94504 148792 94556 148844
rect 99472 148792 99524 148844
rect 127992 148860 128044 148912
rect 109684 148792 109736 148844
rect 120724 148792 120776 148844
rect 127072 148792 127124 148844
rect 156052 148860 156104 148912
rect 165988 148860 166040 148912
rect 177304 148860 177356 148912
rect 183652 148860 183704 148912
rect 211712 148860 211764 148912
rect 222016 148860 222068 148912
rect 232504 148860 232556 148912
rect 238852 148860 238904 148912
rect 268016 148860 268068 148912
rect 277676 148860 277728 148912
rect 289084 148860 289136 148912
rect 306012 148860 306064 148912
rect 316684 148860 316736 148912
rect 323032 148860 323084 148912
rect 352012 148860 352064 148912
rect 361672 148860 361724 148912
rect 373264 148860 373316 148912
rect 379612 148860 379664 148912
rect 408040 148860 408092 148912
rect 417700 148860 417752 148912
rect 428556 148860 428608 148912
rect 434812 148860 434864 148912
rect 463700 148860 463752 148912
rect 474004 148860 474056 148912
rect 485044 148860 485096 148912
rect 501696 148860 501748 148912
rect 512644 148860 512696 148912
rect 518992 148860 519044 148912
rect 547880 148860 547932 148912
rect 137652 148792 137704 148844
rect 148324 148792 148376 148844
rect 193680 148792 193732 148844
rect 204904 148792 204956 148844
rect 249708 148792 249760 148844
rect 260104 148792 260156 148844
rect 333704 148792 333756 148844
rect 344284 148792 344336 148844
rect 390008 148792 390060 148844
rect 400864 148792 400916 148844
rect 445668 148792 445720 148844
rect 456064 148792 456116 148844
rect 529664 148792 529716 148844
rect 540244 148792 540296 148844
rect 36728 148724 36780 148776
rect 557540 148724 557592 148776
rect 16028 146888 16080 146940
rect 547880 146888 547932 146940
rect 25688 146480 25740 146532
rect 71044 146480 71096 146532
rect 212356 146480 212408 146532
rect 232688 146480 232740 146532
rect 296352 146480 296404 146532
rect 316776 146480 316828 146532
rect 408040 146480 408092 146532
rect 428648 146480 428700 146532
rect 492036 146480 492088 146532
rect 512736 146480 512788 146532
rect 36912 146412 36964 146464
rect 53656 146412 53708 146464
rect 148416 146412 148468 146464
rect 165712 146412 165764 146464
rect 175464 146412 175516 146464
rect 193680 146412 193732 146464
rect 203524 146412 203576 146464
rect 221372 146412 221424 146464
rect 260104 146412 260156 146464
rect 277676 146412 277728 146464
rect 287520 146412 287572 146464
rect 305368 146412 305420 146464
rect 345664 146412 345716 146464
rect 361672 146412 361724 146464
rect 371516 146412 371568 146464
rect 389364 146412 389416 146464
rect 399484 146412 399536 146464
rect 417700 146412 417752 146464
rect 456064 146412 456116 146464
rect 473360 146412 473412 146464
rect 483480 146412 483532 146464
rect 501696 146412 501748 146464
rect 37004 146344 37056 146396
rect 63316 146344 63368 146396
rect 64328 146344 64380 146396
rect 81440 146344 81492 146396
rect 91468 146344 91520 146396
rect 109684 146344 109736 146396
rect 119436 146344 119488 146396
rect 137652 146344 137704 146396
rect 156328 146344 156380 146396
rect 178684 146344 178736 146396
rect 232504 146344 232556 146396
rect 249708 146344 249760 146396
rect 268016 146344 268068 146396
rect 287704 146344 287756 146396
rect 315488 146344 315540 146396
rect 333704 146344 333756 146396
rect 352012 146344 352064 146396
rect 374644 146344 374696 146396
rect 428464 146344 428516 146396
rect 445668 146344 445720 146396
rect 464344 146344 464396 146396
rect 483664 146344 483716 146396
rect 511448 146344 511500 146396
rect 529664 146344 529716 146396
rect 543004 146344 543056 146396
rect 557540 146344 557592 146396
rect 69664 146276 69716 146328
rect 91100 146276 91152 146328
rect 94504 146276 94556 146328
rect 119344 146276 119396 146328
rect 120724 146276 120776 146328
rect 147312 146276 147364 146328
rect 148324 146276 148376 146328
rect 175372 146276 175424 146328
rect 177304 146276 177356 146328
rect 203340 146276 203392 146328
rect 204904 146276 204956 146328
rect 231032 146276 231084 146328
rect 232596 146276 232648 146328
rect 259368 146276 259420 146328
rect 260196 146276 260248 146328
rect 287336 146276 287388 146328
rect 289084 146276 289136 146328
rect 315028 146276 315080 146328
rect 316684 146276 316736 146328
rect 343364 146276 343416 146328
rect 344284 146276 344336 146328
rect 371332 146276 371384 146328
rect 373264 146276 373316 146328
rect 399024 146276 399076 146328
rect 400864 146276 400916 146328
rect 427360 146276 427412 146328
rect 428556 146276 428608 146328
rect 455328 146276 455380 146328
rect 456156 146276 456208 146328
rect 483020 146276 483072 146328
rect 485044 146276 485096 146328
rect 511356 146276 511408 146328
rect 512644 146276 512696 146328
rect 539324 146276 539376 146328
rect 540244 146276 540296 146328
rect 567200 146276 567252 146328
rect 37924 144168 37976 144220
rect 545764 144168 545816 144220
rect 35624 143556 35676 143608
rect 36728 143556 36780 143608
rect 63592 128256 63644 128308
rect 64328 128256 64380 128308
rect 147680 128256 147732 128308
rect 148416 128256 148468 128308
rect 232688 126896 232740 126948
rect 239772 126896 239824 126948
rect 483664 126896 483716 126948
rect 491668 126896 491720 126948
rect 512736 126896 512788 126948
rect 519636 126896 519688 126948
rect 428648 126216 428700 126268
rect 435732 126216 435784 126268
rect 287704 126080 287756 126132
rect 295708 126080 295760 126132
rect 316776 126080 316828 126132
rect 323676 126080 323728 126132
rect 13728 125536 13780 125588
rect 66260 125536 66312 125588
rect 70308 125536 70360 125588
rect 121460 125536 121512 125588
rect 126888 125536 126940 125588
rect 178040 125536 178092 125588
rect 209688 125536 209740 125588
rect 262220 125536 262272 125588
rect 266268 125536 266320 125588
rect 317420 125536 317472 125588
rect 322848 125536 322900 125588
rect 374000 125536 374052 125588
rect 405648 125536 405700 125588
rect 458180 125536 458232 125588
rect 489828 125536 489880 125588
rect 542360 125536 542412 125588
rect 42708 125468 42760 125520
rect 93860 125468 93912 125520
rect 97908 125468 97960 125520
rect 149060 125468 149112 125520
rect 154488 125468 154540 125520
rect 205640 125468 205692 125520
rect 238668 125468 238720 125520
rect 289820 125468 289872 125520
rect 293868 125468 293920 125520
rect 345020 125468 345072 125520
rect 350448 125468 350500 125520
rect 401600 125468 401652 125520
rect 434628 125468 434680 125520
rect 485780 125468 485832 125520
rect 518808 125468 518860 125520
rect 569960 125468 570012 125520
rect 182088 125400 182140 125452
rect 233240 125400 233292 125452
rect 378048 125400 378100 125452
rect 429200 125400 429252 125452
rect 462228 125400 462280 125452
rect 513380 125400 513432 125452
rect 35624 124788 35676 124840
rect 36912 124788 36964 124840
rect 343548 124788 343600 124840
rect 345664 124788 345716 124840
rect 178684 122748 178736 122800
rect 184020 122748 184072 122800
rect 231584 122748 231636 122800
rect 232504 122748 232556 122800
rect 374644 122748 374696 122800
rect 379704 122748 379756 122800
rect 539324 122748 539376 122800
rect 543004 122748 543056 122800
rect 36820 122680 36872 122732
rect 557540 122680 557592 122732
rect 15200 122612 15252 122664
rect 43996 122612 44048 122664
rect 25688 122544 25740 122596
rect 37004 122544 37056 122596
rect 42892 122544 42944 122596
rect 53656 122544 53708 122596
rect 69664 122544 69716 122596
rect 71872 122612 71924 122664
rect 100024 122612 100076 122664
rect 71964 122544 72016 122596
rect 81992 122544 82044 122596
rect 94504 122544 94556 122596
rect 99472 122544 99524 122596
rect 127992 122612 128044 122664
rect 109684 122544 109736 122596
rect 120724 122544 120776 122596
rect 127072 122544 127124 122596
rect 155960 122612 156012 122664
rect 165988 122612 166040 122664
rect 177304 122612 177356 122664
rect 183652 122612 183704 122664
rect 211712 122612 211764 122664
rect 221924 122612 221976 122664
rect 232596 122612 232648 122664
rect 238852 122612 238904 122664
rect 268016 122612 268068 122664
rect 277676 122612 277728 122664
rect 289084 122612 289136 122664
rect 306012 122612 306064 122664
rect 316684 122612 316736 122664
rect 323032 122612 323084 122664
rect 352012 122612 352064 122664
rect 361672 122612 361724 122664
rect 373264 122612 373316 122664
rect 379612 122612 379664 122664
rect 408040 122612 408092 122664
rect 417700 122612 417752 122664
rect 428556 122612 428608 122664
rect 434812 122612 434864 122664
rect 463792 122612 463844 122664
rect 474004 122612 474056 122664
rect 485044 122612 485096 122664
rect 501696 122612 501748 122664
rect 512644 122612 512696 122664
rect 518992 122612 519044 122664
rect 547880 122612 547932 122664
rect 137652 122544 137704 122596
rect 148324 122544 148376 122596
rect 193680 122544 193732 122596
rect 204904 122544 204956 122596
rect 249708 122544 249760 122596
rect 260196 122544 260248 122596
rect 333704 122544 333756 122596
rect 344284 122544 344336 122596
rect 390008 122544 390060 122596
rect 400864 122544 400916 122596
rect 445668 122544 445720 122596
rect 456156 122544 456208 122596
rect 529664 122544 529716 122596
rect 540244 122544 540296 122596
rect 39304 122476 39356 122528
rect 567200 122476 567252 122528
rect 16028 119348 16080 119400
rect 547880 119348 547932 119400
rect 25688 118940 25740 118992
rect 261484 118940 261536 118992
rect 148324 118872 148376 118924
rect 165712 118872 165764 118924
rect 175464 118872 175516 118924
rect 193680 118872 193732 118924
rect 203524 118872 203576 118924
rect 221372 118872 221424 118924
rect 408040 118872 408092 118924
rect 428648 118872 428700 118924
rect 492036 118872 492088 118924
rect 512736 118872 512788 118924
rect 36912 118804 36964 118856
rect 53656 118804 53708 118856
rect 64328 118804 64380 118856
rect 81440 118804 81492 118856
rect 91468 118804 91520 118856
rect 109684 118804 109736 118856
rect 119436 118804 119488 118856
rect 137652 118804 137704 118856
rect 156328 118804 156380 118856
rect 178684 118804 178736 118856
rect 232596 118804 232648 118856
rect 249708 118804 249760 118856
rect 260104 118804 260156 118856
rect 277676 118804 277728 118856
rect 287520 118804 287572 118856
rect 305368 118804 305420 118856
rect 315488 118804 315540 118856
rect 333704 118804 333756 118856
rect 345664 118804 345716 118856
rect 361672 118804 361724 118856
rect 371516 118804 371568 118856
rect 389364 118804 389416 118856
rect 399484 118804 399536 118856
rect 417700 118804 417752 118856
rect 456156 118804 456208 118856
rect 473360 118804 473412 118856
rect 483480 118804 483532 118856
rect 501696 118804 501748 118856
rect 37004 118736 37056 118788
rect 63316 118736 63368 118788
rect 66904 118736 66956 118788
rect 91100 118736 91152 118788
rect 94504 118736 94556 118788
rect 119344 118736 119396 118788
rect 120724 118736 120776 118788
rect 147312 118736 147364 118788
rect 148416 118736 148468 118788
rect 175372 118736 175424 118788
rect 177304 118736 177356 118788
rect 203340 118736 203392 118788
rect 204904 118736 204956 118788
rect 231032 118736 231084 118788
rect 232504 118736 232556 118788
rect 259368 118736 259420 118788
rect 268016 118736 268068 118788
rect 287704 118736 287756 118788
rect 296352 118736 296404 118788
rect 316776 118736 316828 118788
rect 352012 118736 352064 118788
rect 374644 118736 374696 118788
rect 428464 118736 428516 118788
rect 445668 118736 445720 118788
rect 464344 118736 464396 118788
rect 483664 118736 483716 118788
rect 511448 118736 511500 118788
rect 529664 118736 529716 118788
rect 543004 118736 543056 118788
rect 557540 118736 557592 118788
rect 212356 118668 212408 118720
rect 232688 118668 232740 118720
rect 260196 118668 260248 118720
rect 287336 118668 287388 118720
rect 289084 118668 289136 118720
rect 315028 118668 315080 118720
rect 316684 118668 316736 118720
rect 343364 118668 343416 118720
rect 344284 118668 344336 118720
rect 371332 118668 371384 118720
rect 373264 118668 373316 118720
rect 399024 118668 399076 118720
rect 400864 118668 400916 118720
rect 427360 118668 427412 118720
rect 428556 118668 428608 118720
rect 455328 118668 455380 118720
rect 456064 118668 456116 118720
rect 483020 118668 483072 118720
rect 485044 118668 485096 118720
rect 511356 118668 511408 118720
rect 512644 118668 512696 118720
rect 539324 118668 539376 118720
rect 540244 118668 540296 118720
rect 567200 118668 567252 118720
rect 37924 116560 37976 116612
rect 545764 116560 545816 116612
rect 35624 116084 35676 116136
rect 36820 116084 36872 116136
rect 63592 100240 63644 100292
rect 64328 100240 64380 100292
rect 455696 100240 455748 100292
rect 456156 100240 456208 100292
rect 316776 98880 316828 98932
rect 323676 98880 323728 98932
rect 287704 98744 287756 98796
rect 295708 98744 295760 98796
rect 428648 98608 428700 98660
rect 435732 98608 435784 98660
rect 483664 98608 483716 98660
rect 491668 98608 491720 98660
rect 512736 98540 512788 98592
rect 519636 98540 519688 98592
rect 232688 98200 232740 98252
rect 239772 98200 239824 98252
rect 13728 97928 13780 97980
rect 66260 97928 66312 97980
rect 97908 97928 97960 97980
rect 149060 97928 149112 97980
rect 154488 97928 154540 97980
rect 205640 97928 205692 97980
rect 209688 97928 209740 97980
rect 262220 97928 262272 97980
rect 266268 97928 266320 97980
rect 317420 97928 317472 97980
rect 322848 97928 322900 97980
rect 374000 97928 374052 97980
rect 405648 97928 405700 97980
rect 458180 97928 458232 97980
rect 489828 97928 489880 97980
rect 542360 97928 542412 97980
rect 42708 97860 42760 97912
rect 93860 97860 93912 97912
rect 126888 97860 126940 97912
rect 178040 97860 178092 97912
rect 182088 97860 182140 97912
rect 233240 97860 233292 97912
rect 238668 97860 238720 97912
rect 289820 97860 289872 97912
rect 293868 97860 293920 97912
rect 345020 97860 345072 97912
rect 378048 97860 378100 97912
rect 429200 97860 429252 97912
rect 462228 97860 462280 97912
rect 513380 97860 513432 97912
rect 518808 97860 518860 97912
rect 569960 97860 570012 97912
rect 70308 97792 70360 97844
rect 121460 97792 121512 97844
rect 231676 97792 231728 97844
rect 232596 97792 232648 97844
rect 350448 97792 350500 97844
rect 401600 97792 401652 97844
rect 434628 97792 434680 97844
rect 485780 97792 485832 97844
rect 539508 97792 539560 97844
rect 543004 97792 543056 97844
rect 35624 97656 35676 97708
rect 36912 97656 36964 97708
rect 343640 97656 343692 97708
rect 345664 97656 345716 97708
rect 178684 95140 178736 95192
rect 184020 95140 184072 95192
rect 374644 95140 374696 95192
rect 379704 95140 379756 95192
rect 15200 95072 15252 95124
rect 43996 95072 44048 95124
rect 71044 95072 71096 95124
rect 567200 95072 567252 95124
rect 25688 95004 25740 95056
rect 37004 95004 37056 95056
rect 53656 95004 53708 95056
rect 66904 95004 66956 95056
rect 71872 95004 71924 95056
rect 100024 95004 100076 95056
rect 42892 94936 42944 94988
rect 72056 94936 72108 94988
rect 81992 94936 82044 94988
rect 94504 94936 94556 94988
rect 99472 94936 99524 94988
rect 127992 95004 128044 95056
rect 109684 94936 109736 94988
rect 120724 94936 120776 94988
rect 127072 94936 127124 94988
rect 156052 95004 156104 95056
rect 165988 95004 166040 95056
rect 177304 95004 177356 95056
rect 183652 95004 183704 95056
rect 211712 95004 211764 95056
rect 222016 95004 222068 95056
rect 232504 95004 232556 95056
rect 238852 95004 238904 95056
rect 268016 95004 268068 95056
rect 277676 95004 277728 95056
rect 289084 95004 289136 95056
rect 306012 95004 306064 95056
rect 316684 95004 316736 95056
rect 323032 95004 323084 95056
rect 352012 95004 352064 95056
rect 361672 95004 361724 95056
rect 373264 95004 373316 95056
rect 379612 95004 379664 95056
rect 408040 95004 408092 95056
rect 417700 95004 417752 95056
rect 428556 95004 428608 95056
rect 434812 95004 434864 95056
rect 463700 95004 463752 95056
rect 474004 95004 474056 95056
rect 485044 95004 485096 95056
rect 501696 95004 501748 95056
rect 512644 95004 512696 95056
rect 518992 95004 519044 95056
rect 547880 95004 547932 95056
rect 137652 94936 137704 94988
rect 148416 94936 148468 94988
rect 193680 94936 193732 94988
rect 204904 94936 204956 94988
rect 249708 94936 249760 94988
rect 260196 94936 260248 94988
rect 333704 94936 333756 94988
rect 344284 94936 344336 94988
rect 390008 94936 390060 94988
rect 400864 94936 400916 94988
rect 445668 94936 445720 94988
rect 456064 94936 456116 94988
rect 529664 94936 529716 94988
rect 540244 94936 540296 94988
rect 36728 94868 36780 94920
rect 557540 94868 557592 94920
rect 15292 91740 15344 91792
rect 547880 91740 547932 91792
rect 25688 91264 25740 91316
rect 71044 91264 71096 91316
rect 212356 91264 212408 91316
rect 232688 91264 232740 91316
rect 296352 91264 296404 91316
rect 316776 91264 316828 91316
rect 408040 91264 408092 91316
rect 428648 91264 428700 91316
rect 36912 91196 36964 91248
rect 53656 91196 53708 91248
rect 148324 91196 148376 91248
rect 165712 91196 165764 91248
rect 175464 91196 175516 91248
rect 193680 91196 193732 91248
rect 203524 91196 203576 91248
rect 221372 91196 221424 91248
rect 260196 91196 260248 91248
rect 277676 91196 277728 91248
rect 287520 91196 287572 91248
rect 305368 91196 305420 91248
rect 345664 91196 345716 91248
rect 361672 91196 361724 91248
rect 371516 91196 371568 91248
rect 389364 91196 389416 91248
rect 399484 91196 399536 91248
rect 417700 91196 417752 91248
rect 456156 91196 456208 91248
rect 473360 91196 473412 91248
rect 483480 91196 483532 91248
rect 501696 91196 501748 91248
rect 511448 91196 511500 91248
rect 529664 91196 529716 91248
rect 37004 91128 37056 91180
rect 63316 91128 63368 91180
rect 64328 91128 64380 91180
rect 81440 91128 81492 91180
rect 91468 91128 91520 91180
rect 109684 91128 109736 91180
rect 119436 91128 119488 91180
rect 137652 91128 137704 91180
rect 156328 91128 156380 91180
rect 178684 91128 178736 91180
rect 232596 91128 232648 91180
rect 249708 91128 249760 91180
rect 268016 91128 268068 91180
rect 287704 91128 287756 91180
rect 315488 91128 315540 91180
rect 333704 91128 333756 91180
rect 352012 91128 352064 91180
rect 374644 91128 374696 91180
rect 428464 91128 428516 91180
rect 445668 91128 445720 91180
rect 464344 91128 464396 91180
rect 483664 91128 483716 91180
rect 492036 91128 492088 91180
rect 512736 91128 512788 91180
rect 543004 91128 543056 91180
rect 557540 91128 557592 91180
rect 69664 91060 69716 91112
rect 91100 91060 91152 91112
rect 94504 91060 94556 91112
rect 119344 91060 119396 91112
rect 120724 91060 120776 91112
rect 147312 91060 147364 91112
rect 148416 91060 148468 91112
rect 175372 91060 175424 91112
rect 177304 91060 177356 91112
rect 203340 91060 203392 91112
rect 204904 91060 204956 91112
rect 231032 91060 231084 91112
rect 232504 91060 232556 91112
rect 259368 91060 259420 91112
rect 260104 91060 260156 91112
rect 287336 91060 287388 91112
rect 289084 91060 289136 91112
rect 315028 91060 315080 91112
rect 316684 91060 316736 91112
rect 343364 91060 343416 91112
rect 344284 91060 344336 91112
rect 371332 91060 371384 91112
rect 373264 91060 373316 91112
rect 399024 91060 399076 91112
rect 400864 91060 400916 91112
rect 427360 91060 427412 91112
rect 428556 91060 428608 91112
rect 455328 91060 455380 91112
rect 456064 91060 456116 91112
rect 483020 91060 483072 91112
rect 485044 91060 485096 91112
rect 511356 91060 511408 91112
rect 512644 91060 512696 91112
rect 539324 91060 539376 91112
rect 540244 91060 540296 91112
rect 567200 91060 567252 91112
rect 37924 90312 37976 90364
rect 545764 90312 545816 90364
rect 35624 88408 35676 88460
rect 36728 88408 36780 88460
rect 42708 88408 42760 88460
rect 93860 88408 93912 88460
rect 154488 88408 154540 88460
rect 205640 88408 205692 88460
rect 238668 88408 238720 88460
rect 289820 88408 289872 88460
rect 293868 88408 293920 88460
rect 345020 88408 345072 88460
rect 350448 88408 350500 88460
rect 401600 88408 401652 88460
rect 434628 88408 434680 88460
rect 485780 88408 485832 88460
rect 13728 88340 13780 88392
rect 66260 88340 66312 88392
rect 70308 88340 70360 88392
rect 121460 88340 121512 88392
rect 126888 88340 126940 88392
rect 178040 88340 178092 88392
rect 209688 88340 209740 88392
rect 262220 88340 262272 88392
rect 322848 88340 322900 88392
rect 374000 88340 374052 88392
rect 405648 88340 405700 88392
rect 458180 88340 458232 88392
rect 518808 88340 518860 88392
rect 569960 88340 570012 88392
rect 3148 84192 3200 84244
rect 11796 84192 11848 84244
rect 428648 72428 428700 72480
rect 435732 72428 435784 72480
rect 63592 72292 63644 72344
rect 64328 72292 64380 72344
rect 232688 72292 232740 72344
rect 239772 72292 239824 72344
rect 259736 72292 259788 72344
rect 260196 72292 260248 72344
rect 316776 72292 316828 72344
rect 323676 72292 323728 72344
rect 455696 72292 455748 72344
rect 456156 72292 456208 72344
rect 483664 72224 483716 72276
rect 491668 72224 491720 72276
rect 287704 72088 287756 72140
rect 295708 72088 295760 72140
rect 512736 72088 512788 72140
rect 519636 72088 519688 72140
rect 35624 71680 35676 71732
rect 36912 71680 36964 71732
rect 97908 71680 97960 71732
rect 149060 71680 149112 71732
rect 182088 71680 182140 71732
rect 233240 71680 233292 71732
rect 266268 71680 266320 71732
rect 317420 71680 317472 71732
rect 343548 71680 343600 71732
rect 345664 71680 345716 71732
rect 378048 71680 378100 71732
rect 429200 71680 429252 71732
rect 489828 71680 489880 71732
rect 542360 71680 542412 71732
rect 231676 71612 231728 71664
rect 232596 71612 232648 71664
rect 462228 71612 462280 71664
rect 513380 71612 513432 71664
rect 42892 68960 42944 69012
rect 15200 68892 15252 68944
rect 43996 68892 44048 68944
rect 72056 68960 72108 69012
rect 99472 68960 99524 69012
rect 71872 68892 71924 68944
rect 100024 68892 100076 68944
rect 127072 68960 127124 69012
rect 127992 68892 128044 68944
rect 183652 68960 183704 69012
rect 156052 68892 156104 68944
rect 165988 68892 166040 68944
rect 177304 68892 177356 68944
rect 178684 68892 178736 68944
rect 184020 68892 184072 68944
rect 374644 68960 374696 69012
rect 379704 68960 379756 69012
rect 539324 68960 539376 69012
rect 543004 68960 543056 69012
rect 211712 68892 211764 68944
rect 222016 68892 222068 68944
rect 232504 68892 232556 68944
rect 249708 68892 249760 68944
rect 260104 68892 260156 68944
rect 261484 68892 261536 68944
rect 567200 68892 567252 68944
rect 25688 68824 25740 68876
rect 37004 68824 37056 68876
rect 53656 68824 53708 68876
rect 69664 68824 69716 68876
rect 81992 68824 82044 68876
rect 94504 68824 94556 68876
rect 109684 68824 109736 68876
rect 120724 68824 120776 68876
rect 137652 68824 137704 68876
rect 148416 68824 148468 68876
rect 193680 68824 193732 68876
rect 204904 68824 204956 68876
rect 238852 68824 238904 68876
rect 268016 68824 268068 68876
rect 277676 68824 277728 68876
rect 289084 68824 289136 68876
rect 306012 68824 306064 68876
rect 316684 68824 316736 68876
rect 323032 68824 323084 68876
rect 352012 68824 352064 68876
rect 361672 68824 361724 68876
rect 373264 68824 373316 68876
rect 379612 68824 379664 68876
rect 408040 68824 408092 68876
rect 417700 68824 417752 68876
rect 428556 68824 428608 68876
rect 434812 68824 434864 68876
rect 463700 68824 463752 68876
rect 474004 68824 474056 68876
rect 485044 68824 485096 68876
rect 501696 68824 501748 68876
rect 512644 68824 512696 68876
rect 518992 68824 519044 68876
rect 547880 68824 547932 68876
rect 333704 68756 333756 68808
rect 344284 68756 344336 68808
rect 390008 68756 390060 68808
rect 400864 68756 400916 68808
rect 445668 68756 445720 68808
rect 456064 68756 456116 68808
rect 529664 68756 529716 68808
rect 540244 68756 540296 68808
rect 36820 68688 36872 68740
rect 557540 68688 557592 68740
rect 16028 65492 16080 65544
rect 547880 65492 547932 65544
rect 25688 65152 25740 65204
rect 261484 65152 261536 65204
rect 36912 65084 36964 65136
rect 53656 65084 53708 65136
rect 148416 65084 148468 65136
rect 165620 65084 165672 65136
rect 175464 65084 175516 65136
rect 193680 65084 193732 65136
rect 203524 65084 203576 65136
rect 221372 65084 221424 65136
rect 408040 65084 408092 65136
rect 428648 65084 428700 65136
rect 36820 65016 36872 65068
rect 63316 65016 63368 65068
rect 64420 65016 64472 65068
rect 81440 65016 81492 65068
rect 91468 65016 91520 65068
rect 109684 65016 109736 65068
rect 119436 65016 119488 65068
rect 137652 65016 137704 65068
rect 156328 65016 156380 65068
rect 178684 65016 178736 65068
rect 232504 65016 232556 65068
rect 249708 65016 249760 65068
rect 260104 65016 260156 65068
rect 277676 65016 277728 65068
rect 287520 65016 287572 65068
rect 305368 65016 305420 65068
rect 315488 65016 315540 65068
rect 333704 65016 333756 65068
rect 345664 65016 345716 65068
rect 361672 65016 361724 65068
rect 371516 65016 371568 65068
rect 389364 65016 389416 65068
rect 399484 65016 399536 65068
rect 417700 65016 417752 65068
rect 456156 65016 456208 65068
rect 473544 65016 473596 65068
rect 483480 65016 483532 65068
rect 501696 65016 501748 65068
rect 511448 65016 511500 65068
rect 529664 65016 529716 65068
rect 35348 64948 35400 65000
rect 64328 64948 64380 65000
rect 66904 64948 66956 65000
rect 91100 64948 91152 65000
rect 94504 64948 94556 65000
rect 119344 64948 119396 65000
rect 120724 64948 120776 65000
rect 147312 64948 147364 65000
rect 148324 64948 148376 65000
rect 175280 64948 175332 65000
rect 177304 64948 177356 65000
rect 203340 64948 203392 65000
rect 204904 64948 204956 65000
rect 231032 64948 231084 65000
rect 232596 64948 232648 65000
rect 259368 64948 259420 65000
rect 268016 64948 268068 65000
rect 287704 64948 287756 65000
rect 296352 64948 296404 65000
rect 316776 64948 316828 65000
rect 352012 64948 352064 65000
rect 374644 64948 374696 65000
rect 428464 64948 428516 65000
rect 445668 64948 445720 65000
rect 464344 64948 464396 65000
rect 483664 64948 483716 65000
rect 492036 64948 492088 65000
rect 512736 64948 512788 65000
rect 543004 64948 543056 65000
rect 557540 64948 557592 65000
rect 212264 64880 212316 64932
rect 232688 64880 232740 64932
rect 260196 64880 260248 64932
rect 287336 64880 287388 64932
rect 289084 64880 289136 64932
rect 315028 64880 315080 64932
rect 316684 64880 316736 64932
rect 343364 64880 343416 64932
rect 344284 64880 344336 64932
rect 371332 64880 371384 64932
rect 373264 64880 373316 64932
rect 399024 64880 399076 64932
rect 400864 64880 400916 64932
rect 427360 64880 427412 64932
rect 428556 64880 428608 64932
rect 455328 64880 455380 64932
rect 456064 64880 456116 64932
rect 483204 64880 483256 64932
rect 485044 64880 485096 64932
rect 511356 64880 511408 64932
rect 512644 64880 512696 64932
rect 539324 64880 539376 64932
rect 540244 64880 540296 64932
rect 567200 64880 567252 64932
rect 37924 62772 37976 62824
rect 545764 62772 545816 62824
rect 182088 62160 182140 62212
rect 233240 62160 233292 62212
rect 350448 62160 350500 62212
rect 401600 62160 401652 62212
rect 42708 62092 42760 62144
rect 93860 62092 93912 62144
rect 97908 62092 97960 62144
rect 149060 62092 149112 62144
rect 154488 62092 154540 62144
rect 205640 62092 205692 62144
rect 238668 62092 238720 62144
rect 289820 62092 289872 62144
rect 293868 62092 293920 62144
rect 345020 62092 345072 62144
rect 378048 62092 378100 62144
rect 429200 62092 429252 62144
rect 434628 62092 434680 62144
rect 485780 62092 485832 62144
rect 489828 62092 489880 62144
rect 542360 62092 542412 62144
rect 63592 50328 63644 50380
rect 64420 50328 64472 50380
rect 147680 50328 147732 50380
rect 148416 50328 148468 50380
rect 455696 50328 455748 50380
rect 456156 50328 456208 50380
rect 232688 44888 232740 44940
rect 239772 44888 239824 44940
rect 428648 44820 428700 44872
rect 435732 44820 435784 44872
rect 512736 44684 512788 44736
rect 519636 44684 519688 44736
rect 483664 44616 483716 44668
rect 491668 44616 491720 44668
rect 3240 44480 3292 44532
rect 8944 44480 8996 44532
rect 287704 44276 287756 44328
rect 295708 44276 295760 44328
rect 316776 44276 316828 44328
rect 323676 44276 323728 44328
rect 13728 44072 13780 44124
rect 66260 44072 66312 44124
rect 70308 44072 70360 44124
rect 121460 44072 121512 44124
rect 126888 44072 126940 44124
rect 178040 44072 178092 44124
rect 209688 44072 209740 44124
rect 262220 44072 262272 44124
rect 266268 44072 266320 44124
rect 317420 44072 317472 44124
rect 322848 44072 322900 44124
rect 374000 44072 374052 44124
rect 405648 44072 405700 44124
rect 458180 44072 458232 44124
rect 462228 44072 462280 44124
rect 513380 44072 513432 44124
rect 518808 44072 518860 44124
rect 569960 44072 570012 44124
rect 35624 44004 35676 44056
rect 36912 44004 36964 44056
rect 343548 44004 343600 44056
rect 345664 44004 345716 44056
rect 539508 44004 539560 44056
rect 543004 44004 543056 44056
rect 25688 41352 25740 41404
rect 36820 41352 36872 41404
rect 178684 41352 178736 41404
rect 184020 41352 184072 41404
rect 374644 41352 374696 41404
rect 379704 41352 379756 41404
rect 15200 41284 15252 41336
rect 43996 41284 44048 41336
rect 71044 41284 71096 41336
rect 567200 41284 567252 41336
rect 53656 41216 53708 41268
rect 66904 41216 66956 41268
rect 71872 41216 71924 41268
rect 100024 41216 100076 41268
rect 42892 41148 42944 41200
rect 72056 41148 72108 41200
rect 81992 41148 82044 41200
rect 94504 41148 94556 41200
rect 99472 41148 99524 41200
rect 127992 41216 128044 41268
rect 109684 41148 109736 41200
rect 120724 41148 120776 41200
rect 127072 41148 127124 41200
rect 156052 41216 156104 41268
rect 165988 41216 166040 41268
rect 177304 41216 177356 41268
rect 183652 41216 183704 41268
rect 211712 41216 211764 41268
rect 222016 41216 222068 41268
rect 232596 41216 232648 41268
rect 238852 41216 238904 41268
rect 268016 41216 268068 41268
rect 277676 41216 277728 41268
rect 289084 41216 289136 41268
rect 306012 41216 306064 41268
rect 316684 41216 316736 41268
rect 323032 41216 323084 41268
rect 352012 41216 352064 41268
rect 361672 41216 361724 41268
rect 373264 41216 373316 41268
rect 379612 41216 379664 41268
rect 408040 41216 408092 41268
rect 417700 41216 417752 41268
rect 428556 41216 428608 41268
rect 434812 41216 434864 41268
rect 463700 41216 463752 41268
rect 474004 41216 474056 41268
rect 485044 41216 485096 41268
rect 501696 41216 501748 41268
rect 512644 41216 512696 41268
rect 518992 41216 519044 41268
rect 547880 41216 547932 41268
rect 137652 41148 137704 41200
rect 148324 41148 148376 41200
rect 193680 41148 193732 41200
rect 204904 41148 204956 41200
rect 249708 41148 249760 41200
rect 260196 41148 260248 41200
rect 333704 41148 333756 41200
rect 344284 41148 344336 41200
rect 390008 41148 390060 41200
rect 400864 41148 400916 41200
rect 445668 41148 445720 41200
rect 456064 41148 456116 41200
rect 529664 41148 529716 41200
rect 540244 41148 540296 41200
rect 36728 41080 36780 41132
rect 557540 41080 557592 41132
rect 21180 38360 21232 38412
rect 36544 38360 36596 38412
rect 11796 38292 11848 38344
rect 34060 38292 34112 38344
rect 40040 38292 40092 38344
rect 60740 38292 60792 38344
rect 13084 38224 13136 38276
rect 52736 38224 52788 38276
rect 3424 38156 3476 38208
rect 49516 38156 49568 38208
rect 3516 38088 3568 38140
rect 59176 38088 59228 38140
rect 6184 38020 6236 38072
rect 17960 38020 18012 38072
rect 24400 38020 24452 38072
rect 234620 38020 234672 38072
rect 3700 37952 3752 38004
rect 37280 37952 37332 38004
rect 46296 37952 46348 38004
rect 567844 37952 567896 38004
rect 16028 37884 16080 37936
rect 547972 37884 548024 37936
rect 212356 37476 212408 37528
rect 232688 37476 232740 37528
rect 408040 37476 408092 37528
rect 428648 37476 428700 37528
rect 30840 37408 30892 37460
rect 36636 37408 36688 37460
rect 148324 37408 148376 37460
rect 165712 37408 165764 37460
rect 175464 37408 175516 37460
rect 193680 37408 193732 37460
rect 203524 37408 203576 37460
rect 221372 37408 221424 37460
rect 260196 37408 260248 37460
rect 277676 37408 277728 37460
rect 287520 37408 287572 37460
rect 305368 37408 305420 37460
rect 345664 37408 345716 37460
rect 361672 37408 361724 37460
rect 371516 37408 371568 37460
rect 389364 37408 389416 37460
rect 399484 37408 399536 37460
rect 417700 37408 417752 37460
rect 456064 37408 456116 37460
rect 473360 37408 473412 37460
rect 483480 37408 483532 37460
rect 501696 37408 501748 37460
rect 27620 37340 27672 37392
rect 62764 37340 62816 37392
rect 64420 37340 64472 37392
rect 81440 37340 81492 37392
rect 91468 37340 91520 37392
rect 109684 37340 109736 37392
rect 126244 37340 126296 37392
rect 137652 37340 137704 37392
rect 156328 37340 156380 37392
rect 178684 37340 178736 37392
rect 232596 37340 232648 37392
rect 249708 37340 249760 37392
rect 268016 37340 268068 37392
rect 287704 37340 287756 37392
rect 296168 37340 296220 37392
rect 316776 37340 316828 37392
rect 322204 37340 322256 37392
rect 333704 37340 333756 37392
rect 352012 37340 352064 37392
rect 374644 37340 374696 37392
rect 428464 37340 428516 37392
rect 445668 37340 445720 37392
rect 464344 37340 464396 37392
rect 483664 37340 483716 37392
rect 492036 37340 492088 37392
rect 512736 37340 512788 37392
rect 518164 37340 518216 37392
rect 529664 37340 529716 37392
rect 543004 37340 543056 37392
rect 557540 37340 557592 37392
rect 1400 37272 1452 37324
rect 39856 37272 39908 37324
rect 43076 37272 43128 37324
rect 91100 37272 91152 37324
rect 93124 37272 93176 37324
rect 119344 37272 119396 37324
rect 120724 37272 120776 37324
rect 147312 37272 147364 37324
rect 148416 37272 148468 37324
rect 175372 37272 175424 37324
rect 177304 37272 177356 37324
rect 203340 37272 203392 37324
rect 204904 37272 204956 37324
rect 231032 37272 231084 37324
rect 232504 37272 232556 37324
rect 259368 37272 259420 37324
rect 260104 37272 260156 37324
rect 287336 37272 287388 37324
rect 289084 37272 289136 37324
rect 315028 37272 315080 37324
rect 316684 37272 316736 37324
rect 343364 37272 343416 37324
rect 344284 37272 344336 37324
rect 371332 37272 371384 37324
rect 373264 37272 373316 37324
rect 399024 37272 399076 37324
rect 400864 37272 400916 37324
rect 427360 37272 427412 37324
rect 428556 37272 428608 37324
rect 455328 37272 455380 37324
rect 456156 37272 456208 37324
rect 483020 37272 483072 37324
rect 485044 37272 485096 37324
rect 511356 37272 511408 37324
rect 512644 37272 512696 37324
rect 539324 37272 539376 37324
rect 547144 37272 547196 37324
rect 567200 37272 567252 37324
rect 3976 36796 4028 36848
rect 63684 36796 63736 36848
rect 3608 36728 3660 36780
rect 63592 36728 63644 36780
rect 3332 36660 3384 36712
rect 63500 36660 63552 36712
rect 37924 36592 37976 36644
rect 545764 36592 545816 36644
rect 13636 36524 13688 36576
rect 580264 36524 580316 36576
rect 3424 36048 3476 36100
rect 61292 36048 61344 36100
rect 13728 35980 13780 36032
rect 93860 35980 93912 36032
rect 20 35912 72 35964
rect 55588 35912 55640 35964
rect 126888 34620 126940 34672
rect 178040 34620 178092 34672
rect 350448 34620 350500 34672
rect 401600 34620 401652 34672
rect 434628 34620 434680 34672
rect 485780 34620 485832 34672
rect 97908 34552 97960 34604
rect 149060 34552 149112 34604
rect 182088 34552 182140 34604
rect 233240 34552 233292 34604
rect 238668 34552 238720 34604
rect 289820 34552 289872 34604
rect 293868 34552 293920 34604
rect 345020 34552 345072 34604
rect 378048 34552 378100 34604
rect 429200 34552 429252 34604
rect 462228 34552 462280 34604
rect 513380 34552 513432 34604
rect 518808 34552 518860 34604
rect 569960 34552 570012 34604
rect 70308 34484 70360 34536
rect 121460 34484 121512 34536
rect 154488 34484 154540 34536
rect 205640 34484 205692 34536
rect 209688 34484 209740 34536
rect 262220 34484 262272 34536
rect 266268 34484 266320 34536
rect 317420 34484 317472 34536
rect 322848 34484 322900 34536
rect 374000 34484 374052 34536
rect 405648 34484 405700 34536
rect 458180 34484 458232 34536
rect 489828 34484 489880 34536
rect 542360 34484 542412 34536
rect 7564 33056 7616 33108
rect 12440 33056 12492 33108
rect 63500 27548 63552 27600
rect 68284 27548 68336 27600
rect 259736 21428 259788 21480
rect 260196 21428 260248 21480
rect 8944 19252 8996 19304
rect 12440 19252 12492 19304
rect 428648 18572 428700 18624
rect 435732 18572 435784 18624
rect 287704 18232 287756 18284
rect 295708 18232 295760 18284
rect 316776 18096 316828 18148
rect 323676 18096 323728 18148
rect 232688 17960 232740 18012
rect 239772 17960 239824 18012
rect 483664 17960 483716 18012
rect 491668 17960 491720 18012
rect 512736 17960 512788 18012
rect 519636 17960 519688 18012
rect 231676 16532 231728 16584
rect 232596 16532 232648 16584
rect 343548 16532 343600 16584
rect 345664 16532 345716 16584
rect 539508 16532 539560 16584
rect 543004 16532 543056 16584
rect 6276 13744 6328 13796
rect 16028 13744 16080 13796
rect 50160 13744 50212 13796
rect 65524 13744 65576 13796
rect 81992 13744 82044 13796
rect 93124 13744 93176 13796
rect 119344 13744 119396 13796
rect 126244 13744 126296 13796
rect 178684 13744 178736 13796
rect 184020 13744 184072 13796
rect 193680 13744 193732 13796
rect 204904 13744 204956 13796
rect 277676 13744 277728 13796
rect 289084 13744 289136 13796
rect 315672 13744 315724 13796
rect 322204 13744 322256 13796
rect 361672 13744 361724 13796
rect 373264 13744 373316 13796
rect 374644 13744 374696 13796
rect 379704 13744 379756 13796
rect 390008 13744 390060 13796
rect 400864 13744 400916 13796
rect 474004 13744 474056 13796
rect 485044 13744 485096 13796
rect 511356 13744 511408 13796
rect 518164 13744 518216 13796
rect 10324 13676 10376 13728
rect 18604 13676 18656 13728
rect 53380 13676 53432 13728
rect 60740 13676 60792 13728
rect 109684 13676 109736 13728
rect 120724 13676 120776 13728
rect 137652 13676 137704 13728
rect 148416 13676 148468 13728
rect 306012 13676 306064 13728
rect 316684 13676 316736 13728
rect 333704 13676 333756 13728
rect 344284 13676 344336 13728
rect 417700 13676 417752 13728
rect 428556 13676 428608 13728
rect 445668 13676 445720 13728
rect 456156 13676 456208 13728
rect 3884 13608 3936 13660
rect 59820 13608 59872 13660
rect 64328 13608 64380 13660
rect 557540 13608 557592 13660
rect 7656 13540 7708 13592
rect 25044 13540 25096 13592
rect 46940 13540 46992 13592
rect 490564 13540 490616 13592
rect 501696 13540 501748 13592
rect 512644 13540 512696 13592
rect 518992 13540 519044 13592
rect 547880 13540 547932 13592
rect 14464 13472 14516 13524
rect 56600 13472 56652 13524
rect 62764 13472 62816 13524
rect 4804 13404 4856 13456
rect 21824 13404 21876 13456
rect 34704 13404 34756 13456
rect 64144 13404 64196 13456
rect 71872 13472 71924 13524
rect 100024 13472 100076 13524
rect 72056 13404 72108 13456
rect 99472 13404 99524 13456
rect 127992 13472 128044 13524
rect 127072 13404 127124 13456
rect 156052 13472 156104 13524
rect 165988 13472 166040 13524
rect 177304 13472 177356 13524
rect 183652 13472 183704 13524
rect 211712 13472 211764 13524
rect 222016 13472 222068 13524
rect 232504 13472 232556 13524
rect 249708 13472 249760 13524
rect 260104 13472 260156 13524
rect 261484 13472 261536 13524
rect 567200 13472 567252 13524
rect 238852 13404 238904 13456
rect 268016 13404 268068 13456
rect 323032 13404 323084 13456
rect 352012 13404 352064 13456
rect 379612 13404 379664 13456
rect 408040 13404 408092 13456
rect 434812 13404 434864 13456
rect 463700 13404 463752 13456
rect 529664 13404 529716 13456
rect 547144 13404 547196 13456
rect 4068 13336 4120 13388
rect 31484 13336 31536 13388
rect 40500 13336 40552 13388
rect 567936 13336 567988 13388
rect 3792 13268 3844 13320
rect 28264 13268 28316 13320
rect 37924 13268 37976 13320
rect 541624 13268 541676 13320
rect 3424 13064 3476 13116
rect 43720 13064 43772 13116
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 36636 700528 36688 700534
rect 36636 700470 36688 700476
rect 36544 700324 36596 700330
rect 36544 700266 36596 700272
rect 25688 686112 25740 686118
rect 25688 686054 25740 686060
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 25700 683876 25728 686054
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3148 632120 3200 632126
rect 3146 632088 3148 632097
rect 3200 632088 3202 632097
rect 3146 632023 3202 632032
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3252 579766 3280 579935
rect 3240 579760 3292 579766
rect 3240 579702 3292 579708
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3054 306232 3110 306241
rect 3054 306167 3110 306176
rect 3068 305046 3096 306167
rect 3056 305040 3108 305046
rect 3056 304982 3108 304988
rect 3330 254144 3386 254153
rect 3330 254079 3332 254088
rect 3384 254079 3386 254088
rect 3332 254050 3384 254056
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240242 3096 241023
rect 3056 240236 3108 240242
rect 3056 240178 3108 240184
rect 2962 188864 3018 188873
rect 2962 188799 3018 188808
rect 2976 187746 3004 188799
rect 2964 187740 3016 187746
rect 2964 187682 3016 187688
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3238 45520 3294 45529
rect 3238 45455 3294 45464
rect 3252 44538 3280 45455
rect 3240 44532 3292 44538
rect 3240 44474 3292 44480
rect 1400 37324 1452 37330
rect 1400 37266 1452 37272
rect 20 35964 72 35970
rect 20 35906 72 35912
rect 32 16574 60 35906
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 37266
rect 3344 36718 3372 58511
rect 3436 38214 3464 527847
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3424 38208 3476 38214
rect 3424 38150 3476 38156
rect 3528 38146 3556 475623
rect 3606 345400 3662 345409
rect 3606 345335 3662 345344
rect 3516 38140 3568 38146
rect 3516 38082 3568 38088
rect 3620 36786 3648 345335
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3712 38010 3740 293111
rect 3790 201920 3846 201929
rect 3790 201855 3846 201864
rect 3700 38004 3752 38010
rect 3700 37946 3752 37952
rect 3608 36780 3660 36786
rect 3608 36722 3660 36728
rect 3332 36712 3384 36718
rect 3332 36654 3384 36660
rect 3424 36100 3476 36106
rect 3424 36042 3476 36048
rect 3436 19417 3464 36042
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3804 13326 3832 201855
rect 3882 149832 3938 149841
rect 3882 149767 3938 149776
rect 3896 13666 3924 149767
rect 3974 136776 4030 136785
rect 3974 136711 4030 136720
rect 3988 36854 4016 136711
rect 4066 97608 4122 97617
rect 4066 97543 4122 97552
rect 3976 36848 4028 36854
rect 3976 36790 4028 36796
rect 3884 13660 3936 13666
rect 3884 13602 3936 13608
rect 4080 13394 4108 97543
rect 4816 13462 4844 683674
rect 15212 683318 16054 683346
rect 35374 683318 35664 683346
rect 13726 674248 13782 674257
rect 13726 674183 13782 674192
rect 13740 665174 13768 674183
rect 13728 665168 13780 665174
rect 13728 665110 13780 665116
rect 15212 662250 15240 683318
rect 35636 683194 35664 683318
rect 35624 683188 35676 683194
rect 35624 683130 35676 683136
rect 35624 665100 35676 665106
rect 35624 665042 35676 665048
rect 35636 664714 35664 665042
rect 35374 664686 35664 664714
rect 15200 662244 15252 662250
rect 15200 662186 15252 662192
rect 16040 658986 16068 664020
rect 25700 662318 25728 664020
rect 25688 662312 25740 662318
rect 25688 662254 25740 662260
rect 16028 658980 16080 658986
rect 16028 658922 16080 658928
rect 25688 658504 25740 658510
rect 25688 658446 25740 658452
rect 25700 656948 25728 658446
rect 35374 656946 35664 656962
rect 35374 656940 35676 656946
rect 35374 656934 35624 656940
rect 35624 656882 35676 656888
rect 15212 656254 16054 656282
rect 13728 655580 13780 655586
rect 13728 655522 13780 655528
rect 13740 647329 13768 655522
rect 13726 647320 13782 647329
rect 13726 647255 13782 647264
rect 15212 634710 15240 656254
rect 35624 637560 35676 637566
rect 35374 637508 35624 637514
rect 35374 637502 35676 637508
rect 35374 637486 35664 637502
rect 15200 634704 15252 634710
rect 15200 634646 15252 634652
rect 16040 632738 16068 637092
rect 25700 634778 25728 637092
rect 25688 634772 25740 634778
rect 25688 634714 25740 634720
rect 16028 632732 16080 632738
rect 16028 632674 16080 632680
rect 25688 632324 25740 632330
rect 25688 632266 25740 632272
rect 6184 632120 6236 632126
rect 6184 632062 6236 632068
rect 6196 38078 6224 632062
rect 25700 629884 25728 632266
rect 15212 629326 16054 629354
rect 35374 629338 35664 629354
rect 35374 629332 35676 629338
rect 35374 629326 35624 629332
rect 13726 620256 13782 620265
rect 13726 620191 13782 620200
rect 13740 611318 13768 620191
rect 13728 611312 13780 611318
rect 13728 611254 13780 611260
rect 15212 608530 15240 629326
rect 35624 629274 35676 629280
rect 35624 611244 35676 611250
rect 35624 611186 35676 611192
rect 35636 610722 35664 611186
rect 35374 610694 35664 610722
rect 15304 610014 16054 610042
rect 15200 608524 15252 608530
rect 15200 608466 15252 608472
rect 15304 605130 15332 610014
rect 25700 608462 25728 610028
rect 25688 608456 25740 608462
rect 25688 608398 25740 608404
rect 15292 605124 15344 605130
rect 15292 605066 15344 605072
rect 25688 604784 25740 604790
rect 25688 604726 25740 604732
rect 25700 602956 25728 604726
rect 15212 602262 16054 602290
rect 35374 602262 35664 602290
rect 13726 593328 13782 593337
rect 13726 593263 13782 593272
rect 13740 583710 13768 593263
rect 13728 583704 13780 583710
rect 13728 583646 13780 583652
rect 15212 580922 15240 602262
rect 35636 601730 35664 602262
rect 35624 601724 35676 601730
rect 35624 601666 35676 601672
rect 35374 583642 35664 583658
rect 35374 583636 35676 583642
rect 35374 583630 35624 583636
rect 35624 583578 35676 583584
rect 15200 580916 15252 580922
rect 15200 580858 15252 580864
rect 7564 579760 7616 579766
rect 7564 579702 7616 579708
rect 6276 240236 6328 240242
rect 6276 240178 6328 240184
rect 6184 38072 6236 38078
rect 6184 38014 6236 38020
rect 6288 13802 6316 240178
rect 7576 33114 7604 579702
rect 16040 578950 16068 583100
rect 25700 580854 25728 583100
rect 25688 580848 25740 580854
rect 25688 580790 25740 580796
rect 16028 578944 16080 578950
rect 16028 578886 16080 578892
rect 25688 578468 25740 578474
rect 25688 578410 25740 578416
rect 25700 575892 25728 578410
rect 35374 575482 35664 575498
rect 35374 575476 35676 575482
rect 35374 575470 35624 575476
rect 35624 575418 35676 575424
rect 15212 575334 16054 575362
rect 13726 566264 13782 566273
rect 13726 566199 13782 566208
rect 13740 557530 13768 566199
rect 13728 557524 13780 557530
rect 13728 557466 13780 557472
rect 15212 554674 15240 575334
rect 35624 557456 35676 557462
rect 35624 557398 35676 557404
rect 35636 556730 35664 557398
rect 35374 556702 35664 556730
rect 15200 554668 15252 554674
rect 15200 554610 15252 554616
rect 16040 551342 16068 556036
rect 25700 554606 25728 556036
rect 25688 554600 25740 554606
rect 25688 554542 25740 554548
rect 16028 551336 16080 551342
rect 16028 551278 16080 551284
rect 25688 550928 25740 550934
rect 25688 550870 25740 550876
rect 25700 548964 25728 550870
rect 15212 548270 16054 548298
rect 35374 548270 35664 548298
rect 13726 539336 13782 539345
rect 13726 539271 13782 539280
rect 13740 529922 13768 539271
rect 13728 529916 13780 529922
rect 13728 529858 13780 529864
rect 15212 527066 15240 548270
rect 35636 547942 35664 548270
rect 35624 547936 35676 547942
rect 35624 547878 35676 547884
rect 35624 529848 35676 529854
rect 35624 529790 35676 529796
rect 35636 529666 35664 529790
rect 35374 529638 35664 529666
rect 15200 527060 15252 527066
rect 15200 527002 15252 527008
rect 16040 523734 16068 529108
rect 25700 526998 25728 529108
rect 25688 526992 25740 526998
rect 25688 526934 25740 526940
rect 16028 523728 16080 523734
rect 16028 523670 16080 523676
rect 25688 523252 25740 523258
rect 25688 523194 25740 523200
rect 25700 521900 25728 523194
rect 35374 521762 35664 521778
rect 35374 521756 35676 521762
rect 35374 521750 35624 521756
rect 35624 521698 35676 521704
rect 15212 521206 16054 521234
rect 13728 520328 13780 520334
rect 13728 520270 13780 520276
rect 13740 512281 13768 520270
rect 13726 512272 13782 512281
rect 13726 512207 13782 512216
rect 15212 500886 15240 521206
rect 35374 502314 35664 502330
rect 35374 502308 35676 502314
rect 35374 502302 35624 502308
rect 35624 502250 35676 502256
rect 15200 500880 15252 500886
rect 15200 500822 15252 500828
rect 16040 497486 16068 502044
rect 25700 500818 25728 502044
rect 25688 500812 25740 500818
rect 25688 500754 25740 500760
rect 16028 497480 16080 497486
rect 16028 497422 16080 497428
rect 25688 497140 25740 497146
rect 25688 497082 25740 497088
rect 25700 494972 25728 497082
rect 15212 494278 16054 494306
rect 35374 494278 35664 494306
rect 13726 485344 13782 485353
rect 13726 485279 13782 485288
rect 13740 476066 13768 485279
rect 13728 476060 13780 476066
rect 13728 476002 13780 476008
rect 15212 473278 15240 494278
rect 35636 494086 35664 494278
rect 35624 494080 35676 494086
rect 35624 494022 35676 494028
rect 35624 475992 35676 475998
rect 35624 475934 35676 475940
rect 35636 475674 35664 475934
rect 35374 475646 35664 475674
rect 15304 475102 16054 475130
rect 15200 473272 15252 473278
rect 15200 473214 15252 473220
rect 15304 469878 15332 475102
rect 25700 473210 25728 475116
rect 25688 473204 25740 473210
rect 25688 473146 25740 473152
rect 15292 469872 15344 469878
rect 15292 469814 15344 469820
rect 25688 469464 25740 469470
rect 25688 469406 25740 469412
rect 25700 467908 25728 469406
rect 15212 467214 16054 467242
rect 35374 467214 35664 467242
rect 13728 466472 13780 466478
rect 13728 466414 13780 466420
rect 13740 458289 13768 466414
rect 13726 458280 13782 458289
rect 13726 458215 13782 458224
rect 15212 445670 15240 467214
rect 35636 466546 35664 467214
rect 35624 466540 35676 466546
rect 35624 466482 35676 466488
rect 35624 448520 35676 448526
rect 35374 448468 35624 448474
rect 35374 448462 35676 448468
rect 35374 448446 35664 448462
rect 15200 445664 15252 445670
rect 15200 445606 15252 445612
rect 16040 443698 16068 448052
rect 25700 445602 25728 448052
rect 25688 445596 25740 445602
rect 25688 445538 25740 445544
rect 16028 443692 16080 443698
rect 16028 443634 16080 443640
rect 25688 443216 25740 443222
rect 25688 443158 25740 443164
rect 25700 440980 25728 443158
rect 15212 440286 16054 440314
rect 35374 440298 35664 440314
rect 35374 440292 35676 440298
rect 35374 440286 35624 440292
rect 13726 431352 13782 431361
rect 13726 431287 13782 431296
rect 13740 422278 13768 431287
rect 13728 422272 13780 422278
rect 13728 422214 13780 422220
rect 15212 419422 15240 440286
rect 35624 440234 35676 440240
rect 35624 422204 35676 422210
rect 35624 422146 35676 422152
rect 35636 421682 35664 422146
rect 35374 421654 35664 421682
rect 15200 419416 15252 419422
rect 15200 419358 15252 419364
rect 16040 416090 16068 421124
rect 25700 419354 25728 421124
rect 25688 419348 25740 419354
rect 25688 419290 25740 419296
rect 16028 416084 16080 416090
rect 16028 416026 16080 416032
rect 25688 415744 25740 415750
rect 25688 415686 25740 415692
rect 25700 413916 25728 415686
rect 15212 413222 16054 413250
rect 35374 413222 35664 413250
rect 13084 409896 13136 409902
rect 13084 409838 13136 409844
rect 11704 397520 11756 397526
rect 11704 397462 11756 397468
rect 10324 305040 10376 305046
rect 10324 304982 10376 304988
rect 7656 254108 7708 254114
rect 7656 254050 7708 254056
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 7668 13598 7696 254050
rect 8944 44532 8996 44538
rect 8944 44474 8996 44480
rect 8956 19310 8984 44474
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 10336 13734 10364 304982
rect 11716 35873 11744 397462
rect 11796 84244 11848 84250
rect 11796 84186 11848 84192
rect 11808 38350 11836 84186
rect 11796 38344 11848 38350
rect 11796 38286 11848 38292
rect 13096 38282 13124 409838
rect 13726 404288 13782 404297
rect 13726 404223 13782 404232
rect 13740 394670 13768 404223
rect 13728 394664 13780 394670
rect 13728 394606 13780 394612
rect 15212 391882 15240 413222
rect 35636 412690 35664 413222
rect 35624 412684 35676 412690
rect 35624 412626 35676 412632
rect 35374 394602 35664 394618
rect 35374 394596 35676 394602
rect 35374 394590 35624 394596
rect 35624 394538 35676 394544
rect 15200 391876 15252 391882
rect 15200 391818 15252 391824
rect 16040 389842 16068 394060
rect 25700 391950 25728 394060
rect 25688 391944 25740 391950
rect 25688 391886 25740 391892
rect 16028 389836 16080 389842
rect 16028 389778 16080 389784
rect 25688 389428 25740 389434
rect 25688 389370 25740 389376
rect 25700 386852 25728 389370
rect 35374 386442 35664 386458
rect 35374 386436 35676 386442
rect 35374 386430 35624 386436
rect 35624 386378 35676 386384
rect 15580 386294 16054 386322
rect 13726 376816 13782 376825
rect 13726 376751 13782 376760
rect 13740 368490 13768 376751
rect 15580 373994 15608 386294
rect 15212 373966 15608 373994
rect 13728 368484 13780 368490
rect 13728 368426 13780 368432
rect 15212 365634 15240 373966
rect 15200 365628 15252 365634
rect 15200 365570 15252 365576
rect 16040 362234 16068 367132
rect 25700 365702 25728 367132
rect 35374 367118 35664 367146
rect 35636 367062 35664 367118
rect 35624 367056 35676 367062
rect 35624 366998 35676 367004
rect 25688 365696 25740 365702
rect 25688 365638 25740 365644
rect 16028 362228 16080 362234
rect 16028 362170 16080 362176
rect 25688 361888 25740 361894
rect 25688 361830 25740 361836
rect 25700 359924 25728 361830
rect 15212 359230 16054 359258
rect 35374 359230 35664 359258
rect 14464 357468 14516 357474
rect 14464 357410 14516 357416
rect 13726 350296 13782 350305
rect 13726 350231 13782 350240
rect 13740 340882 13768 350231
rect 13728 340876 13780 340882
rect 13728 340818 13780 340824
rect 13726 322960 13782 322969
rect 13726 322895 13782 322904
rect 13740 314634 13768 322895
rect 13728 314628 13780 314634
rect 13728 314570 13780 314576
rect 13726 296304 13782 296313
rect 13726 296239 13782 296248
rect 13740 287026 13768 296239
rect 13728 287020 13780 287026
rect 13728 286962 13780 286968
rect 13728 277432 13780 277438
rect 13728 277374 13780 277380
rect 13740 269249 13768 277374
rect 13726 269240 13782 269249
rect 13726 269175 13782 269184
rect 13726 242312 13782 242321
rect 13726 242247 13782 242256
rect 13740 233238 13768 242247
rect 13728 233232 13780 233238
rect 13728 233174 13780 233180
rect 13726 215248 13782 215257
rect 13726 215183 13782 215192
rect 13740 205630 13768 215183
rect 13728 205624 13780 205630
rect 13728 205566 13780 205572
rect 13726 188320 13782 188329
rect 13726 188255 13782 188264
rect 13176 187740 13228 187746
rect 13176 187682 13228 187688
rect 13084 38276 13136 38282
rect 13084 38218 13136 38224
rect 11702 35864 11758 35873
rect 11702 35799 11758 35808
rect 12440 33108 12492 33114
rect 12440 33050 12492 33056
rect 12452 32473 12480 33050
rect 12438 32464 12494 32473
rect 12438 32399 12494 32408
rect 13188 22273 13216 187682
rect 13740 179382 13768 188255
rect 13728 179376 13780 179382
rect 13728 179318 13780 179324
rect 13726 161256 13782 161265
rect 13726 161191 13782 161200
rect 13740 151774 13768 161191
rect 13728 151768 13780 151774
rect 13728 151710 13780 151716
rect 13726 134328 13782 134337
rect 13726 134263 13782 134272
rect 13740 125594 13768 134263
rect 13728 125588 13780 125594
rect 13728 125530 13780 125536
rect 13726 107264 13782 107273
rect 13726 107199 13782 107208
rect 13740 97986 13768 107199
rect 13728 97980 13780 97986
rect 13728 97922 13780 97928
rect 13728 88392 13780 88398
rect 13728 88334 13780 88340
rect 13740 80345 13768 88334
rect 13726 80336 13782 80345
rect 13726 80271 13782 80280
rect 13726 53272 13782 53281
rect 13726 53207 13782 53216
rect 13740 44130 13768 53207
rect 13728 44124 13780 44130
rect 13728 44066 13780 44072
rect 13636 36576 13688 36582
rect 13636 36518 13688 36524
rect 13648 26234 13676 36518
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13740 29073 13768 35974
rect 13726 29064 13782 29073
rect 13726 28999 13782 29008
rect 13648 26206 13768 26234
rect 13740 25673 13768 26206
rect 13726 25664 13782 25673
rect 13726 25599 13782 25608
rect 13174 22264 13230 22273
rect 13174 22199 13230 22208
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12452 18873 12480 19246
rect 12438 18864 12494 18873
rect 12438 18799 12494 18808
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 7656 13592 7708 13598
rect 7656 13534 7708 13540
rect 14476 13530 14504 357410
rect 15212 338026 15240 359230
rect 35636 358834 35664 359230
rect 35624 358828 35676 358834
rect 35624 358770 35676 358776
rect 35624 340808 35676 340814
rect 35374 340756 35624 340762
rect 35374 340750 35676 340756
rect 35374 340734 35664 340750
rect 15200 338020 15252 338026
rect 15200 337962 15252 337968
rect 16040 336054 16068 340068
rect 25700 337958 25728 340068
rect 25688 337952 25740 337958
rect 25688 337894 25740 337900
rect 16028 336048 16080 336054
rect 16028 335990 16080 335996
rect 25688 335572 25740 335578
rect 25688 335514 25740 335520
rect 25700 332860 25728 335514
rect 35374 332586 35664 332602
rect 35374 332580 35676 332586
rect 35374 332574 35624 332580
rect 35624 332522 35676 332528
rect 15212 332302 16054 332330
rect 15212 311778 15240 332302
rect 35624 314560 35676 314566
rect 35624 314502 35676 314508
rect 35636 313698 35664 314502
rect 35374 313670 35664 313698
rect 15200 311772 15252 311778
rect 15200 311714 15252 311720
rect 16040 308446 16068 313140
rect 25700 311846 25728 313140
rect 25688 311840 25740 311846
rect 25688 311782 25740 311788
rect 16028 308440 16080 308446
rect 16028 308382 16080 308388
rect 25688 308100 25740 308106
rect 25688 308042 25740 308048
rect 25700 305932 25728 308042
rect 15212 305238 16054 305266
rect 35374 305238 35664 305266
rect 15212 284238 15240 305238
rect 35636 305046 35664 305238
rect 35624 305040 35676 305046
rect 35624 304982 35676 304988
rect 35624 286952 35676 286958
rect 35624 286894 35676 286900
rect 35636 286770 35664 286894
rect 35374 286742 35664 286770
rect 15200 284232 15252 284238
rect 15200 284174 15252 284180
rect 16040 280838 16068 286076
rect 25700 284306 25728 286076
rect 25688 284300 25740 284306
rect 25688 284242 25740 284248
rect 16028 280832 16080 280838
rect 16028 280774 16080 280780
rect 25688 280424 25740 280430
rect 25688 280366 25740 280372
rect 25700 278868 25728 280366
rect 15212 278310 16054 278338
rect 35374 278310 35664 278338
rect 15212 256630 15240 278310
rect 35636 277506 35664 278310
rect 35624 277500 35676 277506
rect 35624 277442 35676 277448
rect 35374 259418 35664 259434
rect 35374 259412 35676 259418
rect 35374 259406 35624 259412
rect 35624 259354 35676 259360
rect 15200 256624 15252 256630
rect 15200 256566 15252 256572
rect 16040 254590 16068 259148
rect 25700 256562 25728 259148
rect 25688 256556 25740 256562
rect 25688 256498 25740 256504
rect 16028 254584 16080 254590
rect 16028 254526 16080 254532
rect 25688 254176 25740 254182
rect 25688 254118 25740 254124
rect 25700 251940 25728 254118
rect 15212 251246 16054 251274
rect 35374 251258 35664 251274
rect 35374 251252 35676 251258
rect 35374 251246 35624 251252
rect 15212 230382 15240 251246
rect 35624 251194 35676 251200
rect 35374 232762 35664 232778
rect 35374 232756 35676 232762
rect 35374 232750 35624 232756
rect 35624 232698 35676 232704
rect 15304 232070 16054 232098
rect 15200 230376 15252 230382
rect 15200 230318 15252 230324
rect 15304 227050 15332 232070
rect 25700 230314 25728 232084
rect 25688 230308 25740 230314
rect 25688 230250 25740 230256
rect 15292 227044 15344 227050
rect 15292 226986 15344 226992
rect 25688 226636 25740 226642
rect 25688 226578 25740 226584
rect 25700 224876 25728 226578
rect 15212 224318 16054 224346
rect 35374 224318 35664 224346
rect 15212 202774 15240 224318
rect 35636 223650 35664 224318
rect 35624 223644 35676 223650
rect 35624 223586 35676 223592
rect 35374 205562 35664 205578
rect 35374 205556 35676 205562
rect 35374 205550 35624 205556
rect 35624 205498 35676 205504
rect 15200 202768 15252 202774
rect 15200 202710 15252 202716
rect 16040 200802 16068 205020
rect 25700 202706 25728 205020
rect 25688 202700 25740 202706
rect 25688 202642 25740 202648
rect 16028 200796 16080 200802
rect 16028 200738 16080 200744
rect 25688 200388 25740 200394
rect 25688 200330 25740 200336
rect 25700 197948 25728 200330
rect 35374 197402 35664 197418
rect 35374 197396 35676 197402
rect 35374 197390 35624 197396
rect 35624 197338 35676 197344
rect 15212 197254 16054 197282
rect 15212 176594 15240 197254
rect 35624 179308 35676 179314
rect 35624 179250 35676 179256
rect 35636 178786 35664 179250
rect 35374 178758 35664 178786
rect 15200 176588 15252 176594
rect 15200 176530 15252 176536
rect 16040 173194 16068 178092
rect 25700 176526 25728 178092
rect 25688 176520 25740 176526
rect 25688 176462 25740 176468
rect 16028 173188 16080 173194
rect 16028 173130 16080 173136
rect 25688 172712 25740 172718
rect 25688 172654 25740 172660
rect 25700 170884 25728 172654
rect 15212 170326 16054 170354
rect 35374 170326 35664 170354
rect 15212 148986 15240 170326
rect 35636 169794 35664 170326
rect 35624 169788 35676 169794
rect 35624 169730 35676 169736
rect 35374 151706 35664 151722
rect 35374 151700 35676 151706
rect 35374 151694 35624 151700
rect 35624 151642 35676 151648
rect 15200 148980 15252 148986
rect 15200 148922 15252 148928
rect 16040 146946 16068 151028
rect 25700 148918 25728 151028
rect 25688 148912 25740 148918
rect 25688 148854 25740 148860
rect 16028 146940 16080 146946
rect 16028 146882 16080 146888
rect 25688 146532 25740 146538
rect 25688 146474 25740 146480
rect 25700 143956 25728 146474
rect 35624 143608 35676 143614
rect 35374 143556 35624 143562
rect 35374 143550 35676 143556
rect 35374 143534 35664 143550
rect 15212 143262 16054 143290
rect 15212 122670 15240 143262
rect 35624 124840 35676 124846
rect 35374 124788 35624 124794
rect 35374 124782 35676 124788
rect 35374 124766 35664 124782
rect 15200 122664 15252 122670
rect 15200 122606 15252 122612
rect 16040 119406 16068 124100
rect 25700 122602 25728 124100
rect 25688 122596 25740 122602
rect 25688 122538 25740 122544
rect 16028 119400 16080 119406
rect 16028 119342 16080 119348
rect 25688 118992 25740 118998
rect 25688 118934 25740 118940
rect 25700 116892 25728 118934
rect 15212 116334 16054 116362
rect 35374 116334 35664 116362
rect 15212 95130 15240 116334
rect 35636 116142 35664 116334
rect 35624 116136 35676 116142
rect 35624 116078 35676 116084
rect 35374 97714 35664 97730
rect 35374 97708 35676 97714
rect 35374 97702 35624 97708
rect 35624 97650 35676 97656
rect 15304 97022 16054 97050
rect 15200 95124 15252 95130
rect 15200 95066 15252 95072
rect 15304 91798 15332 97022
rect 25700 95062 25728 97036
rect 25688 95056 25740 95062
rect 25688 94998 25740 95004
rect 15292 91792 15344 91798
rect 15292 91734 15344 91740
rect 25688 91316 25740 91322
rect 25688 91258 25740 91264
rect 25700 89964 25728 91258
rect 15212 89270 16054 89298
rect 35374 89270 35664 89298
rect 15212 68950 15240 89270
rect 35636 88466 35664 89270
rect 35624 88460 35676 88466
rect 35624 88402 35676 88408
rect 35624 71732 35676 71738
rect 35624 71674 35676 71680
rect 35636 70666 35664 71674
rect 35374 70638 35664 70666
rect 15200 68944 15252 68950
rect 15200 68886 15252 68892
rect 16040 65550 16068 70108
rect 25700 68882 25728 70108
rect 25688 68876 25740 68882
rect 25688 68818 25740 68824
rect 16028 65544 16080 65550
rect 16028 65486 16080 65492
rect 25688 65204 25740 65210
rect 25688 65146 25740 65152
rect 25700 62900 25728 65146
rect 35348 65000 35400 65006
rect 35348 64942 35400 64948
rect 35360 62900 35388 64942
rect 15212 62206 16054 62234
rect 15212 41342 15240 62206
rect 35624 44056 35676 44062
rect 35624 43998 35676 44004
rect 35636 43738 35664 43998
rect 35374 43710 35664 43738
rect 15200 41336 15252 41342
rect 15200 41278 15252 41284
rect 16040 37942 16068 43044
rect 25700 41410 25728 43044
rect 25688 41404 25740 41410
rect 25688 41346 25740 41352
rect 36556 38418 36584 700266
rect 21180 38412 21232 38418
rect 21180 38354 21232 38360
rect 36544 38412 36596 38418
rect 36544 38354 36596 38360
rect 17960 38072 18012 38078
rect 17960 38014 18012 38020
rect 16028 37936 16080 37942
rect 16028 37878 16080 37884
rect 17972 35972 18000 38014
rect 21192 35972 21220 38354
rect 34060 38344 34112 38350
rect 34060 38286 34112 38292
rect 24400 38072 24452 38078
rect 24400 38014 24452 38020
rect 24412 35972 24440 38014
rect 30840 37460 30892 37466
rect 30840 37402 30892 37408
rect 27620 37392 27672 37398
rect 27620 37334 27672 37340
rect 27632 35972 27660 37334
rect 30852 35972 30880 37402
rect 34072 35972 34100 38286
rect 36648 37466 36676 700470
rect 36912 686044 36964 686050
rect 36912 685986 36964 685992
rect 36820 685976 36872 685982
rect 36820 685918 36872 685924
rect 36728 683188 36780 683194
rect 36728 683130 36780 683136
rect 36740 634506 36768 683130
rect 36832 662318 36860 685918
rect 36924 665106 36952 685986
rect 37922 673568 37978 673577
rect 37922 673503 37978 673512
rect 36912 665100 36964 665106
rect 36912 665042 36964 665048
rect 36820 662312 36872 662318
rect 36820 662254 36872 662260
rect 37004 658436 37056 658442
rect 37004 658378 37056 658384
rect 36912 658368 36964 658374
rect 36912 658310 36964 658316
rect 36820 656940 36872 656946
rect 36820 656882 36872 656888
rect 36728 634500 36780 634506
rect 36728 634442 36780 634448
rect 36728 629332 36780 629338
rect 36728 629274 36780 629280
rect 36740 580718 36768 629274
rect 36832 608326 36860 656882
rect 36924 634778 36952 658310
rect 37016 637566 37044 658378
rect 37936 657558 37964 673503
rect 37924 657552 37976 657558
rect 37924 657494 37976 657500
rect 37922 646640 37978 646649
rect 37922 646575 37978 646584
rect 37004 637560 37056 637566
rect 37004 637502 37056 637508
rect 36912 634772 36964 634778
rect 36912 634714 36964 634720
rect 37004 632256 37056 632262
rect 37004 632198 37056 632204
rect 36912 632188 36964 632194
rect 36912 632130 36964 632136
rect 36924 608462 36952 632130
rect 37016 611250 37044 632198
rect 37936 629950 37964 646575
rect 37924 629944 37976 629950
rect 37924 629886 37976 629892
rect 37922 619576 37978 619585
rect 37922 619511 37978 619520
rect 37004 611244 37056 611250
rect 37004 611186 37056 611192
rect 36912 608456 36964 608462
rect 36912 608398 36964 608404
rect 36820 608320 36872 608326
rect 36820 608262 36872 608268
rect 37004 604648 37056 604654
rect 37004 604590 37056 604596
rect 36912 604580 36964 604586
rect 36912 604522 36964 604528
rect 36820 601724 36872 601730
rect 36820 601666 36872 601672
rect 36728 580712 36780 580718
rect 36728 580654 36780 580660
rect 36728 575476 36780 575482
rect 36728 575418 36780 575424
rect 36740 526862 36768 575418
rect 36832 554470 36860 601666
rect 36924 580854 36952 604522
rect 37016 583642 37044 604590
rect 37936 602410 37964 619511
rect 37924 602404 37976 602410
rect 37924 602346 37976 602352
rect 37922 592648 37978 592657
rect 37922 592583 37978 592592
rect 37004 583636 37056 583642
rect 37004 583578 37056 583584
rect 36912 580848 36964 580854
rect 36912 580790 36964 580796
rect 36912 578400 36964 578406
rect 36912 578342 36964 578348
rect 36924 557462 36952 578342
rect 37004 578332 37056 578338
rect 37004 578274 37056 578280
rect 36912 557456 36964 557462
rect 36912 557398 36964 557404
rect 37016 554606 37044 578274
rect 37936 576162 37964 592583
rect 37924 576156 37976 576162
rect 37924 576098 37976 576104
rect 37922 565584 37978 565593
rect 37922 565519 37978 565528
rect 37004 554600 37056 554606
rect 37004 554542 37056 554548
rect 36820 554464 36872 554470
rect 36820 554406 36872 554412
rect 36820 550792 36872 550798
rect 36820 550734 36872 550740
rect 36832 529854 36860 550734
rect 37004 550724 37056 550730
rect 37004 550666 37056 550672
rect 36912 547936 36964 547942
rect 36912 547878 36964 547884
rect 36820 529848 36872 529854
rect 36820 529790 36872 529796
rect 36728 526856 36780 526862
rect 36728 526798 36780 526804
rect 36728 523184 36780 523190
rect 36728 523126 36780 523132
rect 36740 502314 36768 523126
rect 36820 521756 36872 521762
rect 36820 521698 36872 521704
rect 36728 502308 36780 502314
rect 36728 502250 36780 502256
rect 36728 494080 36780 494086
rect 36728 494022 36780 494028
rect 36740 445466 36768 494022
rect 36832 473074 36860 521698
rect 36924 500682 36952 547878
rect 37016 526998 37044 550666
rect 37936 548554 37964 565519
rect 37924 548548 37976 548554
rect 37924 548490 37976 548496
rect 37922 538656 37978 538665
rect 37922 538591 37978 538600
rect 37004 526992 37056 526998
rect 37004 526934 37056 526940
rect 37004 523116 37056 523122
rect 37004 523058 37056 523064
rect 37016 500818 37044 523058
rect 37936 522306 37964 538591
rect 37924 522300 37976 522306
rect 37924 522242 37976 522248
rect 37922 511592 37978 511601
rect 37922 511527 37978 511536
rect 37004 500812 37056 500818
rect 37004 500754 37056 500760
rect 36912 500676 36964 500682
rect 36912 500618 36964 500624
rect 37004 497004 37056 497010
rect 37004 496946 37056 496952
rect 36912 496936 36964 496942
rect 36912 496878 36964 496884
rect 36924 473210 36952 496878
rect 37016 475998 37044 496946
rect 37936 494766 37964 511527
rect 37924 494760 37976 494766
rect 37924 494702 37976 494708
rect 37922 484664 37978 484673
rect 37922 484599 37978 484608
rect 37004 475992 37056 475998
rect 37004 475934 37056 475940
rect 36912 473204 36964 473210
rect 36912 473146 36964 473152
rect 36820 473068 36872 473074
rect 36820 473010 36872 473016
rect 37004 469396 37056 469402
rect 37004 469338 37056 469344
rect 36912 469328 36964 469334
rect 36912 469270 36964 469276
rect 36820 466540 36872 466546
rect 36820 466482 36872 466488
rect 36728 445460 36780 445466
rect 36728 445402 36780 445408
rect 36728 440292 36780 440298
rect 36728 440234 36780 440240
rect 36740 391678 36768 440234
rect 36832 419218 36860 466482
rect 36924 445602 36952 469270
rect 37016 448526 37044 469338
rect 37936 468518 37964 484599
rect 37924 468512 37976 468518
rect 37924 468454 37976 468460
rect 37922 457600 37978 457609
rect 37922 457535 37978 457544
rect 37004 448520 37056 448526
rect 37004 448462 37056 448468
rect 36912 445596 36964 445602
rect 36912 445538 36964 445544
rect 36912 443148 36964 443154
rect 36912 443090 36964 443096
rect 36924 422210 36952 443090
rect 37004 443080 37056 443086
rect 37004 443022 37056 443028
rect 36912 422204 36964 422210
rect 36912 422146 36964 422152
rect 37016 419354 37044 443022
rect 37936 440910 37964 457535
rect 37924 440904 37976 440910
rect 37924 440846 37976 440852
rect 37922 430672 37978 430681
rect 37922 430607 37978 430616
rect 37004 419348 37056 419354
rect 37004 419290 37056 419296
rect 36820 419212 36872 419218
rect 36820 419154 36872 419160
rect 37004 415608 37056 415614
rect 37004 415550 37056 415556
rect 36912 415540 36964 415546
rect 36912 415482 36964 415488
rect 36820 412684 36872 412690
rect 36820 412626 36872 412632
rect 36728 391672 36780 391678
rect 36728 391614 36780 391620
rect 36728 386436 36780 386442
rect 36728 386378 36780 386384
rect 36740 337822 36768 386378
rect 36832 365430 36860 412626
rect 36924 391950 36952 415482
rect 37016 394602 37044 415550
rect 37936 414730 37964 430607
rect 37924 414724 37976 414730
rect 37924 414666 37976 414672
rect 37922 403608 37978 403617
rect 37922 403543 37978 403552
rect 37004 394596 37056 394602
rect 37004 394538 37056 394544
rect 36912 391944 36964 391950
rect 36912 391886 36964 391892
rect 37004 389360 37056 389366
rect 37004 389302 37056 389308
rect 36912 389292 36964 389298
rect 36912 389234 36964 389240
rect 36924 365702 36952 389234
rect 37016 367062 37044 389302
rect 37936 387122 37964 403543
rect 37924 387116 37976 387122
rect 37924 387058 37976 387064
rect 37922 376000 37978 376009
rect 37922 375935 37978 375944
rect 37004 367056 37056 367062
rect 37004 366998 37056 367004
rect 36912 365696 36964 365702
rect 36912 365638 36964 365644
rect 36820 365424 36872 365430
rect 36820 365366 36872 365372
rect 37004 361752 37056 361758
rect 37004 361694 37056 361700
rect 36820 361684 36872 361690
rect 36820 361626 36872 361632
rect 36832 337958 36860 361626
rect 36912 358828 36964 358834
rect 36912 358770 36964 358776
rect 36820 337952 36872 337958
rect 36820 337894 36872 337900
rect 36728 337816 36780 337822
rect 36728 337758 36780 337764
rect 36728 335436 36780 335442
rect 36728 335378 36780 335384
rect 36740 311846 36768 335378
rect 36820 332580 36872 332586
rect 36820 332522 36872 332528
rect 36728 311840 36780 311846
rect 36728 311782 36780 311788
rect 36728 305040 36780 305046
rect 36728 304982 36780 304988
rect 36740 256426 36768 304982
rect 36832 284034 36860 332522
rect 36924 311574 36952 358770
rect 37016 340814 37044 361694
rect 37936 359514 37964 375935
rect 37924 359508 37976 359514
rect 37924 359450 37976 359456
rect 37922 349616 37978 349625
rect 37922 349551 37978 349560
rect 37004 340808 37056 340814
rect 37004 340750 37056 340756
rect 37004 335504 37056 335510
rect 37004 335446 37056 335452
rect 37016 314566 37044 335446
rect 37936 333266 37964 349551
rect 37924 333260 37976 333266
rect 37924 333202 37976 333208
rect 37922 322008 37978 322017
rect 37922 321943 37978 321952
rect 37004 314560 37056 314566
rect 37004 314502 37056 314508
rect 36912 311568 36964 311574
rect 36912 311510 36964 311516
rect 37004 307964 37056 307970
rect 37004 307906 37056 307912
rect 36912 307896 36964 307902
rect 36912 307838 36964 307844
rect 36924 284306 36952 307838
rect 37016 286958 37044 307906
rect 37936 305658 37964 321943
rect 37924 305652 37976 305658
rect 37924 305594 37976 305600
rect 37922 295624 37978 295633
rect 37922 295559 37978 295568
rect 37004 286952 37056 286958
rect 37004 286894 37056 286900
rect 36912 284300 36964 284306
rect 36912 284242 36964 284248
rect 36820 284028 36872 284034
rect 36820 283970 36872 283976
rect 37004 280356 37056 280362
rect 37004 280298 37056 280304
rect 36912 280288 36964 280294
rect 36912 280230 36964 280236
rect 36820 277500 36872 277506
rect 36820 277442 36872 277448
rect 36728 256420 36780 256426
rect 36728 256362 36780 256368
rect 36728 251252 36780 251258
rect 36728 251194 36780 251200
rect 36740 202570 36768 251194
rect 36832 230178 36860 277442
rect 36924 256562 36952 280230
rect 37016 259418 37044 280298
rect 37936 279478 37964 295559
rect 37924 279472 37976 279478
rect 37924 279414 37976 279420
rect 37922 268560 37978 268569
rect 37922 268495 37978 268504
rect 37004 259412 37056 259418
rect 37004 259354 37056 259360
rect 36912 256556 36964 256562
rect 36912 256498 36964 256504
rect 37004 254108 37056 254114
rect 37004 254050 37056 254056
rect 36912 254040 36964 254046
rect 36912 253982 36964 253988
rect 36924 230314 36952 253982
rect 37016 232762 37044 254050
rect 37936 251870 37964 268495
rect 37924 251864 37976 251870
rect 37924 251806 37976 251812
rect 37922 241632 37978 241641
rect 37922 241567 37978 241576
rect 37004 232756 37056 232762
rect 37004 232698 37056 232704
rect 36912 230308 36964 230314
rect 36912 230250 36964 230256
rect 36820 230172 36872 230178
rect 36820 230114 36872 230120
rect 37004 226500 37056 226506
rect 37004 226442 37056 226448
rect 36912 226432 36964 226438
rect 36912 226374 36964 226380
rect 36820 223644 36872 223650
rect 36820 223586 36872 223592
rect 36728 202564 36780 202570
rect 36728 202506 36780 202512
rect 36728 197396 36780 197402
rect 36728 197338 36780 197344
rect 36740 148782 36768 197338
rect 36832 176390 36860 223586
rect 36924 202706 36952 226374
rect 37016 205562 37044 226442
rect 37936 225622 37964 241567
rect 37924 225616 37976 225622
rect 37924 225558 37976 225564
rect 37922 214568 37978 214577
rect 37922 214503 37978 214512
rect 37004 205556 37056 205562
rect 37004 205498 37056 205504
rect 36912 202700 36964 202706
rect 36912 202642 36964 202648
rect 36912 200320 36964 200326
rect 36912 200262 36964 200268
rect 36924 179314 36952 200262
rect 37004 200252 37056 200258
rect 37004 200194 37056 200200
rect 36912 179308 36964 179314
rect 36912 179250 36964 179256
rect 37016 176526 37044 200194
rect 37936 198014 37964 214503
rect 37924 198008 37976 198014
rect 37924 197950 37976 197956
rect 37922 187640 37978 187649
rect 37922 187575 37978 187584
rect 37004 176520 37056 176526
rect 37004 176462 37056 176468
rect 36820 176384 36872 176390
rect 36820 176326 36872 176332
rect 37004 172644 37056 172650
rect 37004 172586 37056 172592
rect 36912 172576 36964 172582
rect 36912 172518 36964 172524
rect 36820 169788 36872 169794
rect 36820 169730 36872 169736
rect 36728 148776 36780 148782
rect 36728 148718 36780 148724
rect 36728 143608 36780 143614
rect 36728 143550 36780 143556
rect 36740 94926 36768 143550
rect 36832 122738 36860 169730
rect 36924 148918 36952 172518
rect 37016 151706 37044 172586
rect 37936 170406 37964 187575
rect 39304 172712 39356 172718
rect 39304 172654 39356 172660
rect 37924 170400 37976 170406
rect 37924 170342 37976 170348
rect 37922 160576 37978 160585
rect 37922 160511 37978 160520
rect 37004 151700 37056 151706
rect 37004 151642 37056 151648
rect 36912 148912 36964 148918
rect 36912 148854 36964 148860
rect 36912 146464 36964 146470
rect 36912 146406 36964 146412
rect 36924 124846 36952 146406
rect 37004 146396 37056 146402
rect 37004 146338 37056 146344
rect 36912 124840 36964 124846
rect 36912 124782 36964 124788
rect 36820 122732 36872 122738
rect 36820 122674 36872 122680
rect 37016 122602 37044 146338
rect 37936 144226 37964 160511
rect 37924 144220 37976 144226
rect 37924 144162 37976 144168
rect 37922 133648 37978 133657
rect 37922 133583 37978 133592
rect 37004 122596 37056 122602
rect 37004 122538 37056 122544
rect 36912 118856 36964 118862
rect 36912 118798 36964 118804
rect 36820 116136 36872 116142
rect 36820 116078 36872 116084
rect 36728 94920 36780 94926
rect 36728 94862 36780 94868
rect 36728 88460 36780 88466
rect 36728 88402 36780 88408
rect 36740 41138 36768 88402
rect 36832 68746 36860 116078
rect 36924 97714 36952 118798
rect 37004 118788 37056 118794
rect 37004 118730 37056 118736
rect 36912 97708 36964 97714
rect 36912 97650 36964 97656
rect 37016 95062 37044 118730
rect 37936 116618 37964 133583
rect 39316 122534 39344 172654
rect 39304 122528 39356 122534
rect 39304 122470 39356 122476
rect 37924 116612 37976 116618
rect 37924 116554 37976 116560
rect 37922 106584 37978 106593
rect 37922 106519 37978 106528
rect 37004 95056 37056 95062
rect 37004 94998 37056 95004
rect 36912 91248 36964 91254
rect 36912 91190 36964 91196
rect 36924 71738 36952 91190
rect 37004 91180 37056 91186
rect 37004 91122 37056 91128
rect 36912 71732 36964 71738
rect 36912 71674 36964 71680
rect 37016 68882 37044 91122
rect 37936 90370 37964 106519
rect 37924 90364 37976 90370
rect 37924 90306 37976 90312
rect 37922 79656 37978 79665
rect 37922 79591 37978 79600
rect 37004 68876 37056 68882
rect 37004 68818 37056 68824
rect 36820 68740 36872 68746
rect 36820 68682 36872 68688
rect 36912 65136 36964 65142
rect 36912 65078 36964 65084
rect 36820 65068 36872 65074
rect 36820 65010 36872 65016
rect 36832 41410 36860 65010
rect 36924 44062 36952 65078
rect 37936 62830 37964 79591
rect 37924 62824 37976 62830
rect 37924 62766 37976 62772
rect 37922 52592 37978 52601
rect 37922 52527 37978 52536
rect 36912 44056 36964 44062
rect 36912 43998 36964 44004
rect 36820 41404 36872 41410
rect 36820 41346 36872 41352
rect 36728 41132 36780 41138
rect 36728 41074 36780 41080
rect 37280 38004 37332 38010
rect 37280 37946 37332 37952
rect 36636 37460 36688 37466
rect 36636 37402 36688 37408
rect 37292 35972 37320 37946
rect 37936 36650 37964 52527
rect 40052 38350 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 105464 700670 105492 703520
rect 68284 700664 68336 700670
rect 68284 700606 68336 700612
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 64144 700596 64196 700602
rect 64144 700538 64196 700544
rect 53656 686044 53708 686050
rect 53656 685986 53708 685992
rect 53668 683876 53696 685986
rect 63316 685976 63368 685982
rect 63316 685918 63368 685924
rect 63328 683876 63356 685918
rect 42904 683318 44022 683346
rect 42708 683188 42760 683194
rect 42708 683130 42760 683136
rect 42720 674257 42748 683130
rect 42706 674248 42762 674257
rect 42706 674183 42762 674192
rect 42904 662318 42932 683318
rect 63592 668772 63644 668778
rect 63592 668714 63644 668720
rect 63604 664714 63632 668714
rect 63342 664686 63632 664714
rect 43640 664006 44022 664034
rect 53576 664006 53682 664034
rect 42892 662312 42944 662318
rect 42892 662254 42944 662260
rect 43640 662250 43668 664006
rect 53576 663794 53604 664006
rect 53576 663766 53788 663794
rect 53760 662318 53788 663766
rect 53748 662312 53800 662318
rect 53748 662254 53800 662260
rect 43628 662244 43680 662250
rect 43628 662186 43680 662192
rect 53656 658436 53708 658442
rect 53656 658378 53708 658384
rect 53668 656948 53696 658378
rect 63316 658368 63368 658374
rect 63316 658310 63368 658316
rect 63328 656948 63356 658310
rect 42904 656254 44022 656282
rect 42708 655648 42760 655654
rect 42708 655590 42760 655596
rect 42720 647329 42748 655590
rect 42706 647320 42762 647329
rect 42706 647255 42762 647264
rect 42904 634574 42932 656254
rect 63592 640824 63644 640830
rect 63592 640766 63644 640772
rect 63604 637786 63632 640766
rect 63342 637758 63632 637786
rect 44008 634710 44036 637092
rect 43996 634704 44048 634710
rect 43996 634646 44048 634652
rect 53668 634642 53696 637092
rect 53656 634636 53708 634642
rect 53656 634578 53708 634584
rect 42892 634568 42944 634574
rect 42892 634510 42944 634516
rect 53656 632256 53708 632262
rect 53656 632198 53708 632204
rect 53668 629884 53696 632198
rect 63316 632188 63368 632194
rect 63316 632130 63368 632136
rect 63328 629884 63356 632130
rect 42904 629326 44022 629354
rect 42706 620256 42762 620265
rect 42706 620191 42762 620200
rect 42720 611250 42748 620191
rect 42708 611244 42760 611250
rect 42708 611186 42760 611192
rect 42904 608462 42932 629326
rect 63592 612808 63644 612814
rect 63592 612750 63644 612756
rect 63604 610722 63632 612750
rect 63342 610694 63632 610722
rect 44008 608530 44036 610028
rect 43996 608524 44048 608530
rect 43996 608466 44048 608472
rect 42892 608456 42944 608462
rect 42892 608398 42944 608404
rect 53668 608394 53696 610028
rect 53656 608388 53708 608394
rect 53656 608330 53708 608336
rect 53656 604648 53708 604654
rect 53656 604590 53708 604596
rect 53668 602956 53696 604590
rect 63316 604580 63368 604586
rect 63316 604522 63368 604528
rect 63328 602956 63356 604522
rect 42904 602262 44022 602290
rect 42706 593328 42762 593337
rect 42706 593263 42762 593272
rect 42720 583642 42748 593263
rect 42708 583636 42760 583642
rect 42708 583578 42760 583584
rect 42904 580786 42932 602262
rect 63592 583704 63644 583710
rect 63342 583652 63592 583658
rect 63342 583646 63644 583652
rect 63342 583630 63632 583646
rect 44008 580922 44036 583100
rect 43996 580916 44048 580922
rect 43996 580858 44048 580864
rect 53668 580854 53696 583100
rect 53656 580848 53708 580854
rect 53656 580790 53708 580796
rect 42892 580780 42944 580786
rect 42892 580722 42944 580728
rect 53656 578400 53708 578406
rect 53656 578342 53708 578348
rect 53668 575892 53696 578342
rect 63316 578332 63368 578338
rect 63316 578274 63368 578280
rect 63328 575892 63356 578274
rect 42904 575334 44022 575362
rect 42706 566264 42762 566273
rect 42706 566199 42762 566208
rect 42720 557462 42748 566199
rect 42708 557456 42760 557462
rect 42708 557398 42760 557404
rect 42904 554742 42932 575334
rect 63592 558340 63644 558346
rect 63592 558282 63644 558288
rect 63604 556730 63632 558282
rect 63342 556702 63632 556730
rect 42892 554736 42944 554742
rect 42892 554678 42944 554684
rect 44008 554674 44036 556036
rect 43996 554668 44048 554674
rect 43996 554610 44048 554616
rect 53668 554606 53696 556036
rect 53656 554600 53708 554606
rect 53656 554542 53708 554548
rect 53656 550792 53708 550798
rect 53656 550734 53708 550740
rect 53668 548964 53696 550734
rect 63316 550724 63368 550730
rect 63316 550666 63368 550672
rect 63328 548964 63356 550666
rect 42904 548270 44022 548298
rect 42706 539336 42762 539345
rect 42706 539271 42762 539280
rect 42720 529854 42748 539271
rect 42708 529848 42760 529854
rect 42708 529790 42760 529796
rect 42904 526930 42932 548270
rect 63592 533656 63644 533662
rect 63592 533598 63644 533604
rect 63604 529666 63632 533598
rect 63342 529638 63632 529666
rect 44008 527066 44036 529108
rect 43996 527060 44048 527066
rect 43996 527002 44048 527008
rect 53668 526998 53696 529108
rect 53656 526992 53708 526998
rect 53656 526934 53708 526940
rect 42892 526924 42944 526930
rect 42892 526866 42944 526872
rect 53656 523184 53708 523190
rect 53656 523126 53708 523132
rect 53668 521900 53696 523126
rect 63316 523116 63368 523122
rect 63316 523058 63368 523064
rect 63328 521900 63356 523058
rect 42904 521206 44022 521234
rect 42708 520396 42760 520402
rect 42708 520338 42760 520344
rect 42720 512281 42748 520338
rect 42706 512272 42762 512281
rect 42706 512207 42762 512216
rect 42904 500954 42932 521206
rect 63592 505640 63644 505646
rect 63592 505582 63644 505588
rect 63604 502738 63632 505582
rect 63342 502710 63632 502738
rect 42892 500948 42944 500954
rect 42892 500890 42944 500896
rect 44008 500886 44036 502044
rect 43996 500880 44048 500886
rect 43996 500822 44048 500828
rect 53668 500818 53696 502044
rect 53656 500812 53708 500818
rect 53656 500754 53708 500760
rect 53656 497004 53708 497010
rect 53656 496946 53708 496952
rect 53668 494972 53696 496946
rect 63316 496936 63368 496942
rect 63316 496878 63368 496884
rect 63328 494972 63356 496878
rect 42904 494278 44022 494306
rect 42706 485344 42762 485353
rect 42706 485279 42762 485288
rect 42720 475998 42748 485279
rect 42708 475992 42760 475998
rect 42708 475934 42760 475940
rect 42904 473142 42932 494278
rect 63592 477692 63644 477698
rect 63592 477634 63644 477640
rect 63604 475674 63632 477634
rect 63342 475646 63632 475674
rect 44008 473278 44036 475116
rect 43996 473272 44048 473278
rect 43996 473214 44048 473220
rect 53668 473210 53696 475116
rect 53656 473204 53708 473210
rect 53656 473146 53708 473152
rect 42892 473136 42944 473142
rect 42892 473078 42944 473084
rect 53656 469396 53708 469402
rect 53656 469338 53708 469344
rect 53668 467908 53696 469338
rect 63316 469328 63368 469334
rect 63316 469270 63368 469276
rect 63328 467908 63356 469270
rect 42904 467214 44022 467242
rect 42708 466540 42760 466546
rect 42708 466482 42760 466488
rect 42720 458289 42748 466482
rect 42706 458280 42762 458289
rect 42706 458215 42762 458224
rect 42904 445738 42932 467214
rect 63592 449676 63644 449682
rect 63592 449618 63644 449624
rect 63604 448746 63632 449618
rect 63342 448718 63632 448746
rect 42892 445732 42944 445738
rect 42892 445674 42944 445680
rect 44008 445670 44036 448052
rect 43996 445664 44048 445670
rect 43996 445606 44048 445612
rect 53668 445602 53696 448052
rect 53656 445596 53708 445602
rect 53656 445538 53708 445544
rect 53380 443148 53432 443154
rect 53380 443090 53432 443096
rect 53392 440994 53420 443090
rect 62948 443080 63000 443086
rect 62948 443022 63000 443028
rect 62960 440994 62988 443022
rect 53392 440966 53682 440994
rect 62960 440966 63342 440994
rect 42708 440292 42760 440298
rect 42708 440234 42760 440240
rect 42904 440286 44022 440314
rect 42720 431361 42748 440234
rect 42706 431352 42762 431361
rect 42706 431287 42762 431296
rect 42904 419286 42932 440286
rect 63592 427168 63644 427174
rect 63592 427110 63644 427116
rect 63604 421682 63632 427110
rect 63342 421654 63632 421682
rect 44008 419422 44036 421124
rect 43996 419416 44048 419422
rect 43996 419358 44048 419364
rect 53668 419354 53696 421124
rect 53656 419348 53708 419354
rect 53656 419290 53708 419296
rect 42892 419280 42944 419286
rect 42892 419222 42944 419228
rect 53656 415608 53708 415614
rect 53656 415550 53708 415556
rect 53668 413916 53696 415550
rect 63316 415540 63368 415546
rect 63316 415482 63368 415488
rect 63328 413916 63356 415482
rect 42904 413222 44022 413250
rect 42706 404288 42762 404297
rect 42706 404223 42762 404232
rect 42720 394602 42748 404223
rect 42708 394596 42760 394602
rect 42708 394538 42760 394544
rect 42904 391746 42932 413222
rect 63592 394664 63644 394670
rect 63342 394612 63592 394618
rect 63342 394606 63644 394612
rect 63342 394590 63632 394606
rect 44008 391882 44036 394060
rect 43996 391876 44048 391882
rect 43996 391818 44048 391824
rect 53668 391814 53696 394060
rect 53656 391808 53708 391814
rect 53656 391750 53708 391756
rect 42892 391740 42944 391746
rect 42892 391682 42944 391688
rect 53656 389360 53708 389366
rect 53656 389302 53708 389308
rect 53668 386852 53696 389302
rect 63316 389292 63368 389298
rect 63316 389234 63368 389240
rect 63328 386852 63356 389234
rect 43548 386294 44022 386322
rect 42706 376816 42762 376825
rect 42706 376751 42762 376760
rect 42720 368422 42748 376751
rect 43548 373994 43576 386294
rect 42904 373966 43576 373994
rect 42708 368416 42760 368422
rect 42708 368358 42760 368364
rect 42904 365702 42932 373966
rect 63592 370592 63644 370598
rect 63592 370534 63644 370540
rect 63604 367690 63632 370534
rect 63342 367662 63632 367690
rect 42892 365696 42944 365702
rect 42892 365638 42944 365644
rect 44008 365634 44036 367132
rect 43996 365628 44048 365634
rect 43996 365570 44048 365576
rect 53668 365566 53696 367132
rect 53656 365560 53708 365566
rect 53656 365502 53708 365508
rect 53656 361752 53708 361758
rect 53656 361694 53708 361700
rect 53668 359924 53696 361694
rect 63316 361684 63368 361690
rect 63316 361626 63368 361632
rect 63328 359924 63356 361626
rect 42904 359230 44022 359258
rect 42706 350296 42762 350305
rect 42706 350231 42762 350240
rect 42720 340814 42748 350231
rect 42708 340808 42760 340814
rect 42708 340750 42760 340756
rect 42904 337890 42932 359230
rect 63592 342576 63644 342582
rect 63592 342518 63644 342524
rect 63604 340762 63632 342518
rect 63342 340734 63632 340762
rect 44008 338026 44036 340068
rect 43996 338020 44048 338026
rect 43996 337962 44048 337968
rect 53668 337958 53696 340068
rect 53656 337952 53708 337958
rect 53656 337894 53708 337900
rect 42892 337884 42944 337890
rect 42892 337826 42944 337832
rect 53656 335504 53708 335510
rect 53656 335446 53708 335452
rect 53668 332860 53696 335446
rect 63316 335436 63368 335442
rect 63316 335378 63368 335384
rect 63328 332860 63356 335378
rect 42904 332302 44022 332330
rect 42706 322960 42762 322969
rect 42706 322895 42762 322904
rect 42720 314566 42748 322895
rect 42708 314560 42760 314566
rect 42708 314502 42760 314508
rect 42904 311846 42932 332302
rect 63592 314696 63644 314702
rect 63592 314638 63644 314644
rect 63604 313698 63632 314638
rect 63342 313670 63632 313698
rect 42892 311840 42944 311846
rect 42892 311782 42944 311788
rect 44008 311778 44036 313140
rect 43996 311772 44048 311778
rect 43996 311714 44048 311720
rect 53668 311710 53696 313140
rect 53656 311704 53708 311710
rect 53656 311646 53708 311652
rect 53656 307964 53708 307970
rect 53656 307906 53708 307912
rect 53668 305932 53696 307906
rect 63316 307896 63368 307902
rect 63316 307838 63368 307844
rect 63328 305932 63356 307838
rect 42904 305238 44022 305266
rect 42706 296304 42762 296313
rect 42706 296239 42762 296248
rect 42720 286958 42748 296239
rect 42708 286952 42760 286958
rect 42708 286894 42760 286900
rect 42904 284102 42932 305238
rect 63592 291916 63644 291922
rect 63592 291858 63644 291864
rect 63604 286770 63632 291858
rect 63342 286742 63632 286770
rect 44008 284238 44036 286076
rect 43996 284232 44048 284238
rect 43996 284174 44048 284180
rect 53668 284170 53696 286076
rect 53656 284164 53708 284170
rect 53656 284106 53708 284112
rect 42892 284096 42944 284102
rect 42892 284038 42944 284044
rect 53656 280356 53708 280362
rect 53656 280298 53708 280304
rect 53668 278868 53696 280298
rect 63316 280288 63368 280294
rect 63316 280230 63368 280236
rect 63328 278868 63356 280230
rect 42904 278310 44022 278338
rect 42708 277500 42760 277506
rect 42708 277442 42760 277448
rect 42720 269249 42748 277442
rect 42706 269240 42762 269249
rect 42706 269175 42762 269184
rect 42904 256698 42932 278310
rect 63592 263492 63644 263498
rect 63592 263434 63644 263440
rect 63604 259706 63632 263434
rect 63342 259678 63632 259706
rect 42892 256692 42944 256698
rect 42892 256634 42944 256640
rect 44008 256630 44036 259148
rect 43996 256624 44048 256630
rect 43996 256566 44048 256572
rect 53668 256562 53696 259148
rect 53656 256556 53708 256562
rect 53656 256498 53708 256504
rect 53656 254108 53708 254114
rect 53656 254050 53708 254056
rect 53668 251940 53696 254050
rect 63316 254040 63368 254046
rect 63316 253982 63368 253988
rect 63328 251940 63356 253982
rect 42708 251252 42760 251258
rect 42708 251194 42760 251200
rect 42904 251246 44022 251274
rect 42720 242321 42748 251194
rect 42706 242312 42762 242321
rect 42706 242247 42762 242256
rect 42904 230246 42932 251246
rect 63592 235408 63644 235414
rect 63592 235350 63644 235356
rect 63604 232778 63632 235350
rect 63342 232750 63632 232778
rect 44008 230382 44036 232084
rect 43996 230376 44048 230382
rect 43996 230318 44048 230324
rect 53668 230314 53696 232084
rect 53656 230308 53708 230314
rect 53656 230250 53708 230256
rect 42892 230240 42944 230246
rect 42892 230182 42944 230188
rect 53656 226500 53708 226506
rect 53656 226442 53708 226448
rect 53668 224876 53696 226442
rect 63316 226432 63368 226438
rect 63316 226374 63368 226380
rect 63328 224876 63356 226374
rect 42904 224318 44022 224346
rect 42706 215248 42762 215257
rect 42706 215183 42762 215192
rect 42720 205562 42748 215183
rect 42708 205556 42760 205562
rect 42708 205498 42760 205504
rect 42904 202638 42932 224318
rect 63592 207392 63644 207398
rect 63592 207334 63644 207340
rect 63604 205578 63632 207334
rect 63342 205550 63632 205578
rect 43640 205006 44022 205034
rect 53576 205006 53682 205034
rect 43640 202774 43668 205006
rect 43628 202768 43680 202774
rect 43628 202710 43680 202716
rect 53576 202706 53604 205006
rect 53564 202700 53616 202706
rect 53564 202642 53616 202648
rect 42892 202632 42944 202638
rect 42892 202574 42944 202580
rect 53656 200320 53708 200326
rect 53656 200262 53708 200268
rect 53668 197948 53696 200262
rect 63316 200252 63368 200258
rect 63316 200194 63368 200200
rect 63328 197948 63356 200194
rect 42904 197254 44022 197282
rect 42706 188320 42762 188329
rect 42706 188255 42762 188264
rect 42720 179314 42748 188255
rect 42708 179308 42760 179314
rect 42708 179250 42760 179256
rect 42904 176662 42932 197254
rect 63592 185632 63644 185638
rect 63592 185574 63644 185580
rect 63604 178786 63632 185574
rect 63342 178758 63632 178786
rect 42892 176656 42944 176662
rect 42892 176598 42944 176604
rect 44008 176594 44036 178092
rect 43996 176588 44048 176594
rect 43996 176530 44048 176536
rect 53668 176526 53696 178092
rect 53656 176520 53708 176526
rect 53656 176462 53708 176468
rect 53656 172644 53708 172650
rect 53656 172586 53708 172592
rect 53668 170884 53696 172586
rect 63316 172576 63368 172582
rect 63316 172518 63368 172524
rect 63328 170884 63356 172518
rect 42904 170326 44022 170354
rect 42706 161256 42762 161265
rect 42706 161191 42762 161200
rect 42720 151706 42748 161191
rect 42708 151700 42760 151706
rect 42708 151642 42760 151648
rect 42904 148850 42932 170326
rect 63592 156664 63644 156670
rect 63592 156606 63644 156612
rect 63604 151722 63632 156606
rect 63342 151694 63632 151722
rect 44008 148986 44036 151028
rect 43996 148980 44048 148986
rect 43996 148922 44048 148928
rect 53668 148918 53696 151028
rect 53656 148912 53708 148918
rect 53656 148854 53708 148860
rect 42892 148844 42944 148850
rect 42892 148786 42944 148792
rect 53656 146464 53708 146470
rect 53656 146406 53708 146412
rect 53668 143956 53696 146406
rect 63316 146396 63368 146402
rect 63316 146338 63368 146344
rect 63328 143956 63356 146338
rect 42904 143262 44022 143290
rect 42706 134328 42762 134337
rect 42706 134263 42762 134272
rect 42720 125526 42748 134263
rect 42708 125520 42760 125526
rect 42708 125462 42760 125468
rect 42904 122602 42932 143262
rect 63592 128308 63644 128314
rect 63592 128250 63644 128256
rect 63604 124794 63632 128250
rect 63342 124766 63632 124794
rect 44008 122670 44036 124100
rect 43996 122664 44048 122670
rect 43996 122606 44048 122612
rect 53668 122602 53696 124100
rect 42892 122596 42944 122602
rect 42892 122538 42944 122544
rect 53656 122596 53708 122602
rect 53656 122538 53708 122544
rect 53656 118856 53708 118862
rect 53656 118798 53708 118804
rect 53668 116892 53696 118798
rect 63316 118788 63368 118794
rect 63316 118730 63368 118736
rect 63328 116892 63356 118730
rect 42904 116334 44022 116362
rect 42706 107264 42762 107273
rect 42706 107199 42762 107208
rect 42720 97918 42748 107199
rect 42708 97912 42760 97918
rect 42708 97854 42760 97860
rect 42904 94994 42932 116334
rect 63592 100292 63644 100298
rect 63592 100234 63644 100240
rect 63604 97730 63632 100234
rect 63342 97702 63632 97730
rect 44008 95130 44036 97036
rect 43996 95124 44048 95130
rect 43996 95066 44048 95072
rect 53668 95062 53696 97036
rect 53656 95056 53708 95062
rect 53656 94998 53708 95004
rect 42892 94988 42944 94994
rect 42892 94930 42944 94936
rect 53656 91248 53708 91254
rect 53656 91190 53708 91196
rect 53668 89964 53696 91190
rect 63316 91180 63368 91186
rect 63316 91122 63368 91128
rect 63328 89964 63356 91122
rect 42904 89270 44022 89298
rect 42708 88460 42760 88466
rect 42708 88402 42760 88408
rect 42720 80345 42748 88402
rect 42706 80336 42762 80345
rect 42706 80271 42762 80280
rect 42904 69018 42932 89270
rect 63592 72344 63644 72350
rect 63592 72286 63644 72292
rect 63604 70666 63632 72286
rect 63342 70638 63632 70666
rect 42892 69012 42944 69018
rect 42892 68954 42944 68960
rect 44008 68950 44036 70108
rect 43996 68944 44048 68950
rect 43996 68886 44048 68892
rect 53668 68882 53696 70108
rect 53656 68876 53708 68882
rect 53656 68818 53708 68824
rect 53656 65136 53708 65142
rect 53656 65078 53708 65084
rect 53668 62900 53696 65078
rect 63316 65068 63368 65074
rect 63316 65010 63368 65016
rect 63328 62900 63356 65010
rect 42904 62206 44022 62234
rect 42708 62144 42760 62150
rect 42708 62086 42760 62092
rect 42720 53281 42748 62086
rect 42706 53272 42762 53281
rect 42706 53207 42762 53216
rect 42904 41206 42932 62206
rect 63592 50380 63644 50386
rect 63592 50322 63644 50328
rect 63604 43738 63632 50322
rect 63342 43710 63632 43738
rect 44008 41342 44036 43044
rect 43996 41336 44048 41342
rect 43996 41278 44048 41284
rect 53668 41274 53696 43044
rect 53656 41268 53708 41274
rect 53656 41210 53708 41216
rect 42892 41200 42944 41206
rect 42892 41142 42944 41148
rect 40040 38344 40092 38350
rect 40040 38286 40092 38292
rect 60740 38344 60792 38350
rect 60740 38286 60792 38292
rect 52736 38276 52788 38282
rect 52736 38218 52788 38224
rect 49516 38208 49568 38214
rect 49516 38150 49568 38156
rect 46296 38004 46348 38010
rect 46296 37946 46348 37952
rect 39856 37324 39908 37330
rect 39856 37266 39908 37272
rect 43076 37324 43128 37330
rect 43076 37266 43128 37272
rect 37924 36644 37976 36650
rect 37924 36586 37976 36592
rect 39868 35972 39896 37266
rect 43088 35972 43116 37266
rect 46308 35972 46336 37946
rect 49528 35972 49556 38150
rect 52748 35972 52776 38218
rect 59176 38140 59228 38146
rect 59176 38082 59228 38088
rect 55600 35970 55982 35986
rect 59188 35972 59216 38082
rect 55588 35964 55982 35970
rect 55640 35958 55982 35964
rect 55588 35906 55640 35912
rect 16040 13802 16068 16116
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 18616 13734 18644 16116
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 21836 13462 21864 16116
rect 25056 13598 25084 16116
rect 25044 13592 25096 13598
rect 25044 13534 25096 13540
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 28276 13326 28304 16116
rect 31496 13394 31524 16116
rect 34716 13462 34744 16116
rect 34704 13456 34756 13462
rect 34704 13398 34756 13404
rect 31484 13388 31536 13394
rect 31484 13330 31536 13336
rect 37936 13326 37964 16116
rect 40512 13394 40540 16116
rect 40500 13388 40552 13394
rect 40500 13330 40552 13336
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 37924 13320 37976 13326
rect 37924 13262 37976 13268
rect 43732 13122 43760 16116
rect 46952 13598 46980 16116
rect 50172 13802 50200 16116
rect 50160 13796 50212 13802
rect 50160 13738 50212 13744
rect 53392 13734 53420 16116
rect 53380 13728 53432 13734
rect 53380 13670 53432 13676
rect 46940 13592 46992 13598
rect 46940 13534 46992 13540
rect 56612 13530 56640 16116
rect 59832 13666 59860 16116
rect 60752 13734 60780 38286
rect 62764 37392 62816 37398
rect 62764 37334 62816 37340
rect 61290 36136 61346 36145
rect 61290 36071 61292 36080
rect 61344 36071 61346 36080
rect 61292 36042 61344 36048
rect 60740 13728 60792 13734
rect 60740 13670 60792 13676
rect 59820 13660 59872 13666
rect 59820 13602 59872 13608
rect 62776 13530 62804 37334
rect 63684 36848 63736 36854
rect 63684 36790 63736 36796
rect 63592 36780 63644 36786
rect 63592 36722 63644 36728
rect 63500 36712 63552 36718
rect 63500 36654 63552 36660
rect 63512 33153 63540 36654
rect 63498 33144 63554 33153
rect 63498 33079 63554 33088
rect 63604 29753 63632 36722
rect 63590 29744 63646 29753
rect 63590 29679 63646 29688
rect 63500 27600 63552 27606
rect 63500 27542 63552 27548
rect 63512 26353 63540 27542
rect 63498 26344 63554 26353
rect 63498 26279 63554 26288
rect 63696 26234 63724 36790
rect 63512 26206 63724 26234
rect 63512 19553 63540 26206
rect 63498 19544 63554 19553
rect 63498 19479 63554 19488
rect 56600 13524 56652 13530
rect 56600 13466 56652 13472
rect 62764 13524 62816 13530
rect 62764 13466 62816 13472
rect 64156 13462 64184 700538
rect 64236 700460 64288 700466
rect 64236 700402 64288 700408
rect 64248 22953 64276 700402
rect 65524 700392 65576 700398
rect 65524 700334 65576 700340
rect 64328 686044 64380 686050
rect 64328 685986 64380 685992
rect 64340 668778 64368 685986
rect 64328 668772 64380 668778
rect 64328 668714 64380 668720
rect 64328 658368 64380 658374
rect 64328 658310 64380 658316
rect 64340 640830 64368 658310
rect 64328 640824 64380 640830
rect 64328 640766 64380 640772
rect 64328 632188 64380 632194
rect 64328 632130 64380 632136
rect 64340 612814 64368 632130
rect 64328 612808 64380 612814
rect 64328 612750 64380 612756
rect 64328 604648 64380 604654
rect 64328 604590 64380 604596
rect 64340 583710 64368 604590
rect 64328 583704 64380 583710
rect 64328 583646 64380 583652
rect 64328 578332 64380 578338
rect 64328 578274 64380 578280
rect 64340 558346 64368 578274
rect 64328 558340 64380 558346
rect 64328 558282 64380 558288
rect 64328 550792 64380 550798
rect 64328 550734 64380 550740
rect 64340 533662 64368 550734
rect 64328 533656 64380 533662
rect 64328 533598 64380 533604
rect 64328 523116 64380 523122
rect 64328 523058 64380 523064
rect 64340 505646 64368 523058
rect 64328 505640 64380 505646
rect 64328 505582 64380 505588
rect 64328 497004 64380 497010
rect 64328 496946 64380 496952
rect 64340 477698 64368 496946
rect 64328 477692 64380 477698
rect 64328 477634 64380 477640
rect 64328 469328 64380 469334
rect 64328 469270 64380 469276
rect 64340 449682 64368 469270
rect 64328 449676 64380 449682
rect 64328 449618 64380 449624
rect 64328 443148 64380 443154
rect 64328 443090 64380 443096
rect 64340 427174 64368 443090
rect 64328 427168 64380 427174
rect 64328 427110 64380 427116
rect 64328 415608 64380 415614
rect 64328 415550 64380 415556
rect 64340 394670 64368 415550
rect 64328 394664 64380 394670
rect 64328 394606 64380 394612
rect 64328 389292 64380 389298
rect 64328 389234 64380 389240
rect 64340 370598 64368 389234
rect 64328 370592 64380 370598
rect 64328 370534 64380 370540
rect 64328 361752 64380 361758
rect 64328 361694 64380 361700
rect 64340 342582 64368 361694
rect 64328 342576 64380 342582
rect 64328 342518 64380 342524
rect 64328 335436 64380 335442
rect 64328 335378 64380 335384
rect 64340 314702 64368 335378
rect 64328 314696 64380 314702
rect 64328 314638 64380 314644
rect 64328 307964 64380 307970
rect 64328 307906 64380 307912
rect 64340 291922 64368 307906
rect 64328 291916 64380 291922
rect 64328 291858 64380 291864
rect 64328 280288 64380 280294
rect 64328 280230 64380 280236
rect 64340 263498 64368 280230
rect 64328 263492 64380 263498
rect 64328 263434 64380 263440
rect 64328 254108 64380 254114
rect 64328 254050 64380 254056
rect 64340 235414 64368 254050
rect 64328 235408 64380 235414
rect 64328 235350 64380 235356
rect 64328 226500 64380 226506
rect 64328 226442 64380 226448
rect 64340 207398 64368 226442
rect 64328 207392 64380 207398
rect 64328 207334 64380 207340
rect 64328 200252 64380 200258
rect 64328 200194 64380 200200
rect 64340 185638 64368 200194
rect 64328 185632 64380 185638
rect 64328 185574 64380 185580
rect 64328 172644 64380 172650
rect 64328 172586 64380 172592
rect 64340 156670 64368 172586
rect 64328 156664 64380 156670
rect 64328 156606 64380 156612
rect 64328 146396 64380 146402
rect 64328 146338 64380 146344
rect 64340 128314 64368 146338
rect 64328 128308 64380 128314
rect 64328 128250 64380 128256
rect 64328 118856 64380 118862
rect 64328 118798 64380 118804
rect 64340 100298 64368 118798
rect 64328 100292 64380 100298
rect 64328 100234 64380 100240
rect 64328 91180 64380 91186
rect 64328 91122 64380 91128
rect 64340 72350 64368 91122
rect 64328 72344 64380 72350
rect 64328 72286 64380 72292
rect 64420 65068 64472 65074
rect 64420 65010 64472 65016
rect 64328 65000 64380 65006
rect 64328 64942 64380 64948
rect 64234 22944 64290 22953
rect 64234 22879 64290 22888
rect 64340 13666 64368 64942
rect 64432 50386 64460 65010
rect 64420 50380 64472 50386
rect 64420 50322 64472 50328
rect 64420 37392 64472 37398
rect 64420 37334 64472 37340
rect 64432 16153 64460 37334
rect 64418 16144 64474 16153
rect 64418 16079 64474 16088
rect 65536 13802 65564 700334
rect 66904 685976 66956 685982
rect 66904 685918 66956 685924
rect 66258 673568 66314 673577
rect 66258 673503 66314 673512
rect 66272 665174 66300 673503
rect 66260 665168 66312 665174
rect 66260 665110 66312 665116
rect 66916 662318 66944 685918
rect 66904 662312 66956 662318
rect 66904 662254 66956 662260
rect 66904 658504 66956 658510
rect 66904 658446 66956 658452
rect 66260 655580 66312 655586
rect 66260 655522 66312 655528
rect 66272 646649 66300 655522
rect 66258 646640 66314 646649
rect 66258 646575 66314 646584
rect 66258 619576 66314 619585
rect 66258 619511 66314 619520
rect 66272 611318 66300 619511
rect 66260 611312 66312 611318
rect 66260 611254 66312 611260
rect 66916 608530 66944 658446
rect 66904 608524 66956 608530
rect 66904 608466 66956 608472
rect 66904 604580 66956 604586
rect 66904 604522 66956 604528
rect 66258 592648 66314 592657
rect 66258 592583 66314 592592
rect 66272 583574 66300 592583
rect 66260 583568 66312 583574
rect 66260 583510 66312 583516
rect 66916 580854 66944 604522
rect 66904 580848 66956 580854
rect 66904 580790 66956 580796
rect 66258 565584 66314 565593
rect 66258 565519 66314 565528
rect 66272 557530 66300 565519
rect 66260 557524 66312 557530
rect 66260 557466 66312 557472
rect 66904 550724 66956 550730
rect 66904 550666 66956 550672
rect 66258 538656 66314 538665
rect 66258 538591 66314 538600
rect 66272 529922 66300 538591
rect 66260 529916 66312 529922
rect 66260 529858 66312 529864
rect 66916 526998 66944 550666
rect 66904 526992 66956 526998
rect 66904 526934 66956 526940
rect 66260 520328 66312 520334
rect 66260 520270 66312 520276
rect 66272 511601 66300 520270
rect 66258 511592 66314 511601
rect 66258 511527 66314 511536
rect 66904 496936 66956 496942
rect 66904 496878 66956 496884
rect 66258 484664 66314 484673
rect 66258 484599 66314 484608
rect 66272 476066 66300 484599
rect 66260 476060 66312 476066
rect 66260 476002 66312 476008
rect 66916 473210 66944 496878
rect 66904 473204 66956 473210
rect 66904 473146 66956 473152
rect 66260 466472 66312 466478
rect 66260 466414 66312 466420
rect 66272 457609 66300 466414
rect 66258 457600 66314 457609
rect 66258 457535 66314 457544
rect 66904 443080 66956 443086
rect 66904 443022 66956 443028
rect 66258 430672 66314 430681
rect 66258 430607 66314 430616
rect 66272 422278 66300 430607
rect 66260 422272 66312 422278
rect 66260 422214 66312 422220
rect 66916 419354 66944 443022
rect 66904 419348 66956 419354
rect 66904 419290 66956 419296
rect 66904 415540 66956 415546
rect 66904 415482 66956 415488
rect 66258 403608 66314 403617
rect 66258 403543 66314 403552
rect 66272 394534 66300 403543
rect 66260 394528 66312 394534
rect 66260 394470 66312 394476
rect 66916 391814 66944 415482
rect 66904 391808 66956 391814
rect 66904 391750 66956 391756
rect 66258 376000 66314 376009
rect 66258 375935 66314 375944
rect 66272 368490 66300 375935
rect 66260 368484 66312 368490
rect 66260 368426 66312 368432
rect 66904 361684 66956 361690
rect 66904 361626 66956 361632
rect 66258 349616 66314 349625
rect 66258 349551 66314 349560
rect 66272 340882 66300 349551
rect 66260 340876 66312 340882
rect 66260 340818 66312 340824
rect 66916 337958 66944 361626
rect 66904 337952 66956 337958
rect 66904 337894 66956 337900
rect 66258 322008 66314 322017
rect 66258 321943 66314 321952
rect 66272 314634 66300 321943
rect 66260 314628 66312 314634
rect 66260 314570 66312 314576
rect 66904 307896 66956 307902
rect 66904 307838 66956 307844
rect 66258 295624 66314 295633
rect 66258 295559 66314 295568
rect 66272 287026 66300 295559
rect 66260 287020 66312 287026
rect 66260 286962 66312 286968
rect 66916 284170 66944 307838
rect 66904 284164 66956 284170
rect 66904 284106 66956 284112
rect 66260 277432 66312 277438
rect 66260 277374 66312 277380
rect 66272 268569 66300 277374
rect 66258 268560 66314 268569
rect 66258 268495 66314 268504
rect 66904 254040 66956 254046
rect 66904 253982 66956 253988
rect 66258 241632 66314 241641
rect 66258 241567 66314 241576
rect 66272 233238 66300 241567
rect 66260 233232 66312 233238
rect 66260 233174 66312 233180
rect 66916 230314 66944 253982
rect 66904 230308 66956 230314
rect 66904 230250 66956 230256
rect 66904 226432 66956 226438
rect 66904 226374 66956 226380
rect 66258 214568 66314 214577
rect 66258 214503 66314 214512
rect 66272 205630 66300 214503
rect 66260 205624 66312 205630
rect 66260 205566 66312 205572
rect 66916 202706 66944 226374
rect 66904 202700 66956 202706
rect 66904 202642 66956 202648
rect 66258 187640 66314 187649
rect 66258 187575 66314 187584
rect 66272 179382 66300 187575
rect 66260 179376 66312 179382
rect 66260 179318 66312 179324
rect 66904 172576 66956 172582
rect 66904 172518 66956 172524
rect 66258 160576 66314 160585
rect 66258 160511 66314 160520
rect 66272 151774 66300 160511
rect 66260 151768 66312 151774
rect 66260 151710 66312 151716
rect 66916 148918 66944 172518
rect 66904 148912 66956 148918
rect 66904 148854 66956 148860
rect 66258 133648 66314 133657
rect 66258 133583 66314 133592
rect 66272 125594 66300 133583
rect 66260 125588 66312 125594
rect 66260 125530 66312 125536
rect 66904 118788 66956 118794
rect 66904 118730 66956 118736
rect 66258 106584 66314 106593
rect 66258 106519 66314 106528
rect 66272 97986 66300 106519
rect 66260 97980 66312 97986
rect 66260 97922 66312 97928
rect 66916 95062 66944 118730
rect 66904 95056 66956 95062
rect 66904 94998 66956 95004
rect 66260 88392 66312 88398
rect 66260 88334 66312 88340
rect 66272 79665 66300 88334
rect 66258 79656 66314 79665
rect 66258 79591 66314 79600
rect 66904 65000 66956 65006
rect 66904 64942 66956 64948
rect 66258 52592 66314 52601
rect 66258 52527 66314 52536
rect 66272 44130 66300 52527
rect 66260 44124 66312 44130
rect 66260 44066 66312 44072
rect 66916 41274 66944 64942
rect 66904 41268 66956 41274
rect 66904 41210 66956 41216
rect 68296 27606 68324 700606
rect 170324 700602 170352 703520
rect 170312 700596 170364 700602
rect 170312 700538 170364 700544
rect 71044 686112 71096 686118
rect 71044 686054 71096 686060
rect 212356 686112 212408 686118
rect 212356 686054 212408 686060
rect 232688 686112 232740 686118
rect 232688 686054 232740 686060
rect 70306 673840 70362 673849
rect 70306 673775 70362 673784
rect 70320 665174 70348 673775
rect 70308 665168 70360 665174
rect 70308 665110 70360 665116
rect 69664 658300 69716 658306
rect 69664 658242 69716 658248
rect 69676 634642 69704 658242
rect 70308 655580 70360 655586
rect 70308 655522 70360 655528
rect 70320 647329 70348 655522
rect 70306 647320 70362 647329
rect 70306 647255 70362 647264
rect 71056 634710 71084 686054
rect 81440 686044 81492 686050
rect 81440 685986 81492 685992
rect 148416 686044 148468 686050
rect 148416 685986 148468 685992
rect 165712 686044 165764 686050
rect 165712 685986 165764 685992
rect 175464 686044 175516 686050
rect 175464 685986 175516 685992
rect 193680 686044 193732 686050
rect 193680 685986 193732 685992
rect 203524 686044 203576 686050
rect 203524 685986 203576 685992
rect 81452 683890 81480 685986
rect 91100 685976 91152 685982
rect 91100 685918 91152 685924
rect 91468 685976 91520 685982
rect 91468 685918 91520 685924
rect 109684 685976 109736 685982
rect 109684 685918 109736 685924
rect 119436 685976 119488 685982
rect 119436 685918 119488 685924
rect 137652 685976 137704 685982
rect 137652 685918 137704 685924
rect 91112 683890 91140 685918
rect 81452 683862 81696 683890
rect 91112 683862 91356 683890
rect 71884 683318 72036 683346
rect 71884 662386 71912 683318
rect 91480 664714 91508 685918
rect 94504 685908 94556 685914
rect 94504 685850 94556 685856
rect 93860 683188 93912 683194
rect 93860 683130 93912 683136
rect 93872 673577 93900 683130
rect 93858 673568 93914 673577
rect 93858 673503 93914 673512
rect 91356 664686 91508 664714
rect 72022 663794 72050 664020
rect 81696 664006 82032 664034
rect 71976 663766 72050 663794
rect 71872 662380 71924 662386
rect 71872 662322 71924 662328
rect 71976 662250 72004 663766
rect 82004 662318 82032 664006
rect 94516 662318 94544 685850
rect 109696 683876 109724 685918
rect 119344 685908 119396 685914
rect 119344 685850 119396 685856
rect 119356 683876 119384 685850
rect 99484 683318 100050 683346
rect 97908 683188 97960 683194
rect 97908 683130 97960 683136
rect 97920 674257 97948 683130
rect 97906 674248 97962 674257
rect 97906 674183 97962 674192
rect 99484 662318 99512 683318
rect 119448 664714 119476 685918
rect 120724 685908 120776 685914
rect 120724 685850 120776 685856
rect 119370 664686 119476 664714
rect 100036 662386 100064 664020
rect 100024 662380 100076 662386
rect 100024 662322 100076 662328
rect 109696 662318 109724 664020
rect 120736 662318 120764 685850
rect 137664 683876 137692 685918
rect 147312 685908 147364 685914
rect 147312 685850 147364 685856
rect 148324 685908 148376 685914
rect 148324 685850 148376 685856
rect 147324 683876 147352 685850
rect 127084 683318 128018 683346
rect 126886 674248 126942 674257
rect 126886 674183 126942 674192
rect 121458 673568 121514 673577
rect 121458 673503 121514 673512
rect 121472 665174 121500 673503
rect 126900 665174 126928 674183
rect 121460 665168 121512 665174
rect 121460 665110 121512 665116
rect 126888 665168 126940 665174
rect 126888 665110 126940 665116
rect 81992 662312 82044 662318
rect 81992 662254 82044 662260
rect 94504 662312 94556 662318
rect 94504 662254 94556 662260
rect 99472 662312 99524 662318
rect 99472 662254 99524 662260
rect 109684 662312 109736 662318
rect 109684 662254 109736 662260
rect 120724 662312 120776 662318
rect 120724 662254 120776 662260
rect 127084 662250 127112 683318
rect 147680 668772 147732 668778
rect 147680 668714 147732 668720
rect 147692 664714 147720 668714
rect 147338 664686 147720 664714
rect 127728 664006 128018 664034
rect 137678 664006 137968 664034
rect 127728 662386 127756 664006
rect 127716 662380 127768 662386
rect 127716 662322 127768 662328
rect 137940 662318 137968 664006
rect 148336 662318 148364 685850
rect 148428 668778 148456 685986
rect 156328 685976 156380 685982
rect 156328 685918 156380 685924
rect 156340 683890 156368 685918
rect 156032 683862 156368 683890
rect 165724 683754 165752 685986
rect 175372 685908 175424 685914
rect 175372 685850 175424 685856
rect 175384 683754 175412 685850
rect 165692 683726 165752 683754
rect 175352 683726 175412 683754
rect 149060 683188 149112 683194
rect 149060 683130 149112 683136
rect 154488 683188 154540 683194
rect 154488 683130 154540 683136
rect 149072 673577 149100 683130
rect 154500 674257 154528 683130
rect 154486 674248 154542 674257
rect 154486 674183 154542 674192
rect 149058 673568 149114 673577
rect 149058 673503 149114 673512
rect 148416 668772 148468 668778
rect 148416 668714 148468 668720
rect 175476 664714 175504 685986
rect 178684 685976 178736 685982
rect 178684 685918 178736 685924
rect 177304 685908 177356 685914
rect 177304 685850 177356 685856
rect 175352 664686 175504 664714
rect 156018 663794 156046 664020
rect 165692 664006 166028 664034
rect 155972 663766 156046 663794
rect 137928 662312 137980 662318
rect 137928 662254 137980 662260
rect 148324 662312 148376 662318
rect 148324 662254 148376 662260
rect 155972 662250 156000 663766
rect 166000 662386 166028 664006
rect 177316 662386 177344 685850
rect 178038 673568 178094 673577
rect 178038 673503 178094 673512
rect 178052 665174 178080 673503
rect 178040 665168 178092 665174
rect 178040 665110 178092 665116
rect 178696 662386 178724 685918
rect 193692 683876 193720 685986
rect 203340 685908 203392 685914
rect 203340 685850 203392 685856
rect 203352 683876 203380 685850
rect 183664 683318 184046 683346
rect 182088 683256 182140 683262
rect 182088 683198 182140 683204
rect 182100 674257 182128 683198
rect 182086 674248 182142 674257
rect 182086 674183 182142 674192
rect 165988 662380 166040 662386
rect 165988 662322 166040 662328
rect 177304 662380 177356 662386
rect 177304 662322 177356 662328
rect 178684 662380 178736 662386
rect 178684 662322 178736 662328
rect 183664 662318 183692 683318
rect 203536 664714 203564 685986
rect 204904 685908 204956 685914
rect 204904 685850 204956 685856
rect 203366 664686 203564 664714
rect 184032 662386 184060 664020
rect 184020 662380 184072 662386
rect 184020 662322 184072 662328
rect 193692 662318 193720 664020
rect 204916 662318 204944 685850
rect 212368 683890 212396 686054
rect 221372 686044 221424 686050
rect 221372 685986 221424 685992
rect 212060 683862 212396 683890
rect 221384 683890 221412 685986
rect 232504 685976 232556 685982
rect 232504 685918 232556 685924
rect 231032 685908 231084 685914
rect 231032 685850 231084 685856
rect 231044 683890 231072 685850
rect 221384 683862 221720 683890
rect 231044 683862 231380 683890
rect 205640 683188 205692 683194
rect 205640 683130 205692 683136
rect 205652 674121 205680 683130
rect 209686 674248 209742 674257
rect 209686 674183 209742 674192
rect 205638 674112 205694 674121
rect 205638 674047 205694 674056
rect 209700 665174 209728 674183
rect 232516 673454 232544 685918
rect 232596 685908 232648 685914
rect 232596 685850 232648 685856
rect 231872 673426 232544 673454
rect 209688 665168 209740 665174
rect 209688 665110 209740 665116
rect 231872 664850 231900 673426
rect 231780 664822 231900 664850
rect 231780 664714 231808 664822
rect 231380 664686 231808 664714
rect 211724 664006 212060 664034
rect 221720 664006 222056 664034
rect 211724 662386 211752 664006
rect 211712 662380 211764 662386
rect 211712 662322 211764 662328
rect 222028 662318 222056 664006
rect 232608 662318 232636 685850
rect 232700 665310 232728 686054
rect 233240 683256 233292 683262
rect 233240 683198 233292 683204
rect 233252 673577 233280 683198
rect 233238 673568 233294 673577
rect 233238 673503 233294 673512
rect 232688 665304 232740 665310
rect 232688 665246 232740 665252
rect 183652 662312 183704 662318
rect 183652 662254 183704 662260
rect 193680 662312 193732 662318
rect 193680 662254 193732 662260
rect 204904 662312 204956 662318
rect 204904 662254 204956 662260
rect 222016 662312 222068 662318
rect 222016 662254 222068 662260
rect 232596 662312 232648 662318
rect 232596 662254 232648 662260
rect 71964 662244 72016 662250
rect 71964 662186 72016 662192
rect 127072 662244 127124 662250
rect 127072 662186 127124 662192
rect 155960 662244 156012 662250
rect 155960 662186 156012 662192
rect 212356 658504 212408 658510
rect 212356 658446 212408 658452
rect 232688 658504 232740 658510
rect 232688 658446 232740 658452
rect 148324 658436 148376 658442
rect 148324 658378 148376 658384
rect 165712 658436 165764 658442
rect 165712 658378 165764 658384
rect 175464 658436 175516 658442
rect 175464 658378 175516 658384
rect 193680 658436 193732 658442
rect 193680 658378 193732 658384
rect 203524 658436 203576 658442
rect 203524 658378 203576 658384
rect 81440 658368 81492 658374
rect 81440 658310 81492 658316
rect 91468 658368 91520 658374
rect 91468 658310 91520 658316
rect 109684 658368 109736 658374
rect 109684 658310 109736 658316
rect 119436 658368 119488 658374
rect 119436 658310 119488 658316
rect 137652 658368 137704 658374
rect 137652 658310 137704 658316
rect 81452 656962 81480 658310
rect 91100 658300 91152 658306
rect 91100 658242 91152 658248
rect 91112 656962 91140 658242
rect 81452 656934 81696 656962
rect 91112 656934 91356 656962
rect 71884 656254 72036 656282
rect 71044 634704 71096 634710
rect 71044 634646 71096 634652
rect 71884 634642 71912 656254
rect 91480 637786 91508 658310
rect 94504 658300 94556 658306
rect 94504 658242 94556 658248
rect 93860 655648 93912 655654
rect 93860 655590 93912 655596
rect 93872 646649 93900 655590
rect 93858 646640 93914 646649
rect 93858 646575 93914 646584
rect 91356 637758 91508 637786
rect 72022 636834 72050 637092
rect 81696 637078 82032 637106
rect 71976 636806 72050 636834
rect 69664 634636 69716 634642
rect 69664 634578 69716 634584
rect 71872 634636 71924 634642
rect 71872 634578 71924 634584
rect 71976 634574 72004 636806
rect 82004 634574 82032 637078
rect 94516 634574 94544 658242
rect 109696 656948 109724 658310
rect 119344 658300 119396 658306
rect 119344 658242 119396 658248
rect 119356 656948 119384 658242
rect 99484 656254 100050 656282
rect 97908 655648 97960 655654
rect 97908 655590 97960 655596
rect 97920 647329 97948 655590
rect 97906 647320 97962 647329
rect 97906 647255 97962 647264
rect 99484 634574 99512 656254
rect 119448 637786 119476 658310
rect 120724 658300 120776 658306
rect 120724 658242 120776 658248
rect 119370 637758 119476 637786
rect 100036 634642 100064 637092
rect 100024 634636 100076 634642
rect 100024 634578 100076 634584
rect 109696 634574 109724 637092
rect 120736 634574 120764 658242
rect 137664 656948 137692 658310
rect 147312 658300 147364 658306
rect 147312 658242 147364 658248
rect 147324 656948 147352 658242
rect 127084 656254 128018 656282
rect 121460 655580 121512 655586
rect 121460 655522 121512 655528
rect 126888 655580 126940 655586
rect 126888 655522 126940 655528
rect 121472 646649 121500 655522
rect 126900 647329 126928 655522
rect 126886 647320 126942 647329
rect 126886 647255 126942 647264
rect 121458 646640 121514 646649
rect 121458 646575 121514 646584
rect 127084 634574 127112 656254
rect 148336 644474 148364 658378
rect 156328 658368 156380 658374
rect 156328 658310 156380 658316
rect 148416 658300 148468 658306
rect 148416 658242 148468 658248
rect 147784 644446 148364 644474
rect 147784 637514 147812 644446
rect 147338 637486 147812 637514
rect 128004 634642 128032 637092
rect 127992 634636 128044 634642
rect 127992 634578 128044 634584
rect 137664 634574 137692 637092
rect 148428 634574 148456 658242
rect 156340 656962 156368 658310
rect 156032 656934 156368 656962
rect 165724 656826 165752 658378
rect 175372 658300 175424 658306
rect 175372 658242 175424 658248
rect 175384 656826 175412 658242
rect 165692 656798 165752 656826
rect 175352 656798 175412 656826
rect 149060 655648 149112 655654
rect 149060 655590 149112 655596
rect 154488 655648 154540 655654
rect 154488 655590 154540 655596
rect 149072 646649 149100 655590
rect 154500 647329 154528 655590
rect 154486 647320 154542 647329
rect 154486 647255 154542 647264
rect 149058 646640 149114 646649
rect 149058 646575 149114 646584
rect 175476 637786 175504 658378
rect 178684 658368 178736 658374
rect 178684 658310 178736 658316
rect 177304 658300 177356 658306
rect 177304 658242 177356 658248
rect 175352 637758 175504 637786
rect 156018 636834 156046 637092
rect 165692 637078 166028 637106
rect 155972 636806 156046 636834
rect 155972 634642 156000 636806
rect 166000 634642 166028 637078
rect 177316 634642 177344 658242
rect 178040 655580 178092 655586
rect 178040 655522 178092 655528
rect 178052 646649 178080 655522
rect 178038 646640 178094 646649
rect 178038 646575 178094 646584
rect 178696 634778 178724 658310
rect 193692 656948 193720 658378
rect 203340 658300 203392 658306
rect 203340 658242 203392 658248
rect 203352 656948 203380 658242
rect 183664 656254 184046 656282
rect 183560 655716 183612 655722
rect 183560 655658 183612 655664
rect 183572 654090 183600 655658
rect 182088 654084 182140 654090
rect 182088 654026 182140 654032
rect 183560 654084 183612 654090
rect 183560 654026 183612 654032
rect 182100 647329 182128 654026
rect 182086 647320 182142 647329
rect 182086 647255 182142 647264
rect 178684 634772 178736 634778
rect 178684 634714 178736 634720
rect 183664 634642 183692 656254
rect 203536 637786 203564 658378
rect 204904 658300 204956 658306
rect 204904 658242 204956 658248
rect 203366 637758 203564 637786
rect 184032 634778 184060 637092
rect 184020 634772 184072 634778
rect 184020 634714 184072 634720
rect 155960 634636 156012 634642
rect 155960 634578 156012 634584
rect 165988 634636 166040 634642
rect 165988 634578 166040 634584
rect 177304 634636 177356 634642
rect 177304 634578 177356 634584
rect 183652 634636 183704 634642
rect 183652 634578 183704 634584
rect 193692 634574 193720 637092
rect 204916 634574 204944 658242
rect 212368 656962 212396 658446
rect 221372 658436 221424 658442
rect 221372 658378 221424 658384
rect 212060 656934 212396 656962
rect 221384 656962 221412 658378
rect 232596 658368 232648 658374
rect 232596 658310 232648 658316
rect 231032 658300 231084 658306
rect 231032 658242 231084 658248
rect 232504 658300 232556 658306
rect 232504 658242 232556 658248
rect 231044 656962 231072 658242
rect 221384 656934 221720 656962
rect 231044 656934 231380 656962
rect 205640 655648 205692 655654
rect 205640 655590 205692 655596
rect 205652 646649 205680 655590
rect 209688 655580 209740 655586
rect 209688 655522 209740 655528
rect 209700 647329 209728 655522
rect 209686 647320 209742 647329
rect 209686 647255 209742 647264
rect 205638 646640 205694 646649
rect 205638 646575 205694 646584
rect 211724 637078 212060 637106
rect 221720 637078 221964 637106
rect 231380 637078 231624 637106
rect 211724 634642 211752 637078
rect 221936 634642 221964 637078
rect 231596 634778 231624 637078
rect 231584 634772 231636 634778
rect 231584 634714 231636 634720
rect 232516 634642 232544 658242
rect 232608 634778 232636 658310
rect 232700 639402 232728 658446
rect 233240 655716 233292 655722
rect 233240 655658 233292 655664
rect 233252 646649 233280 655658
rect 233238 646640 233294 646649
rect 233238 646575 233294 646584
rect 232688 639396 232740 639402
rect 232688 639338 232740 639344
rect 232596 634772 232648 634778
rect 232596 634714 232648 634720
rect 211712 634636 211764 634642
rect 211712 634578 211764 634584
rect 221924 634636 221976 634642
rect 221924 634578 221976 634584
rect 232504 634636 232556 634642
rect 232504 634578 232556 634584
rect 71964 634568 72016 634574
rect 71964 634510 72016 634516
rect 81992 634568 82044 634574
rect 81992 634510 82044 634516
rect 94504 634568 94556 634574
rect 94504 634510 94556 634516
rect 99472 634568 99524 634574
rect 99472 634510 99524 634516
rect 109684 634568 109736 634574
rect 109684 634510 109736 634516
rect 120724 634568 120776 634574
rect 120724 634510 120776 634516
rect 127072 634568 127124 634574
rect 127072 634510 127124 634516
rect 137652 634568 137704 634574
rect 137652 634510 137704 634516
rect 148416 634568 148468 634574
rect 148416 634510 148468 634516
rect 193680 634568 193732 634574
rect 193680 634510 193732 634516
rect 204904 634568 204956 634574
rect 204904 634510 204956 634516
rect 71044 632324 71096 632330
rect 71044 632266 71096 632272
rect 212356 632324 212408 632330
rect 212356 632266 212408 632272
rect 232688 632324 232740 632330
rect 232688 632266 232740 632272
rect 69664 632120 69716 632126
rect 69664 632062 69716 632068
rect 69676 608394 69704 632062
rect 70306 620256 70362 620265
rect 70306 620191 70362 620200
rect 70320 611318 70348 620191
rect 70308 611312 70360 611318
rect 70308 611254 70360 611260
rect 69664 608388 69716 608394
rect 69664 608330 69716 608336
rect 70306 593328 70362 593337
rect 70306 593263 70362 593272
rect 70320 583710 70348 593263
rect 70308 583704 70360 583710
rect 70308 583646 70360 583652
rect 71056 580922 71084 632266
rect 148324 632256 148376 632262
rect 148324 632198 148376 632204
rect 165712 632256 165764 632262
rect 165712 632198 165764 632204
rect 175464 632256 175516 632262
rect 175464 632198 175516 632204
rect 193680 632256 193732 632262
rect 193680 632198 193732 632204
rect 203524 632256 203576 632262
rect 203524 632198 203576 632204
rect 81440 632188 81492 632194
rect 81440 632130 81492 632136
rect 91468 632188 91520 632194
rect 91468 632130 91520 632136
rect 109684 632188 109736 632194
rect 109684 632130 109736 632136
rect 119436 632188 119488 632194
rect 119436 632130 119488 632136
rect 137652 632188 137704 632194
rect 137652 632130 137704 632136
rect 81452 629898 81480 632130
rect 91100 632120 91152 632126
rect 91100 632062 91152 632068
rect 91112 629898 91140 632062
rect 81452 629870 81696 629898
rect 91112 629870 91356 629898
rect 71884 629326 72036 629354
rect 71884 608462 71912 629326
rect 91480 610722 91508 632130
rect 95884 632120 95936 632126
rect 95884 632062 95936 632068
rect 93858 619576 93914 619585
rect 93858 619511 93914 619520
rect 93872 611250 93900 619511
rect 93860 611244 93912 611250
rect 93860 611186 93912 611192
rect 91356 610694 91508 610722
rect 72036 610014 72096 610042
rect 81696 610014 82032 610042
rect 72068 608598 72096 610014
rect 72056 608592 72108 608598
rect 72056 608534 72108 608540
rect 71872 608456 71924 608462
rect 71872 608398 71924 608404
rect 82004 608394 82032 610014
rect 95896 608394 95924 632062
rect 109696 629884 109724 632130
rect 119344 632120 119396 632126
rect 119344 632062 119396 632068
rect 119356 629884 119384 632062
rect 99484 629326 100050 629354
rect 97906 620256 97962 620265
rect 97906 620191 97962 620200
rect 97920 611250 97948 620191
rect 97908 611244 97960 611250
rect 97908 611186 97960 611192
rect 99484 608394 99512 629326
rect 119448 610722 119476 632130
rect 120724 632120 120776 632126
rect 120724 632062 120776 632068
rect 119370 610694 119476 610722
rect 100036 608462 100064 610028
rect 100024 608456 100076 608462
rect 100024 608398 100076 608404
rect 109696 608394 109724 610028
rect 120736 608394 120764 632062
rect 137664 629884 137692 632130
rect 147312 632120 147364 632126
rect 147312 632062 147364 632068
rect 147324 629884 147352 632062
rect 127084 629326 128018 629354
rect 126886 620256 126942 620265
rect 126886 620191 126942 620200
rect 121458 619576 121514 619585
rect 121458 619511 121514 619520
rect 121472 611318 121500 619511
rect 126900 611318 126928 620191
rect 121460 611312 121512 611318
rect 121460 611254 121512 611260
rect 126888 611312 126940 611318
rect 126888 611254 126940 611260
rect 127084 608394 127112 629326
rect 148336 615494 148364 632198
rect 156328 632188 156380 632194
rect 156328 632130 156380 632136
rect 148416 632120 148468 632126
rect 148416 632062 148468 632068
rect 147784 615466 148364 615494
rect 147784 610722 147812 615466
rect 147338 610694 147812 610722
rect 128004 608462 128032 610028
rect 127992 608456 128044 608462
rect 127992 608398 128044 608404
rect 137664 608394 137692 610028
rect 148428 608394 148456 632062
rect 156340 629898 156368 632130
rect 156032 629870 156368 629898
rect 165724 629762 165752 632198
rect 175372 632120 175424 632126
rect 175372 632062 175424 632068
rect 175384 629762 175412 632062
rect 165692 629734 165752 629762
rect 175352 629734 175412 629762
rect 154486 620256 154542 620265
rect 154486 620191 154542 620200
rect 149058 619576 149114 619585
rect 149058 619511 149114 619520
rect 149072 611250 149100 619511
rect 154500 611250 154528 620191
rect 149060 611244 149112 611250
rect 149060 611186 149112 611192
rect 154488 611244 154540 611250
rect 154488 611186 154540 611192
rect 175476 610722 175504 632198
rect 178684 632188 178736 632194
rect 178684 632130 178736 632136
rect 177304 632120 177356 632126
rect 177304 632062 177356 632068
rect 175352 610694 175504 610722
rect 156032 610014 156092 610042
rect 165692 610014 166028 610042
rect 156064 608462 156092 610014
rect 166000 608462 166028 610014
rect 177316 608462 177344 632062
rect 178038 619576 178094 619585
rect 178038 619511 178094 619520
rect 178052 611318 178080 619511
rect 178040 611312 178092 611318
rect 178040 611254 178092 611260
rect 178696 608598 178724 632130
rect 193692 629884 193720 632198
rect 203340 632120 203392 632126
rect 203340 632062 203392 632068
rect 203352 629884 203380 632062
rect 183664 629326 184046 629354
rect 182086 620256 182142 620265
rect 182086 620191 182142 620200
rect 182100 611182 182128 620191
rect 182088 611176 182140 611182
rect 182088 611118 182140 611124
rect 178684 608592 178736 608598
rect 178684 608534 178736 608540
rect 183664 608462 183692 629326
rect 203536 610722 203564 632198
rect 204904 632120 204956 632126
rect 204904 632062 204956 632068
rect 203366 610694 203564 610722
rect 184032 608598 184060 610028
rect 184020 608592 184072 608598
rect 184020 608534 184072 608540
rect 156052 608456 156104 608462
rect 156052 608398 156104 608404
rect 165988 608456 166040 608462
rect 165988 608398 166040 608404
rect 177304 608456 177356 608462
rect 177304 608398 177356 608404
rect 183652 608456 183704 608462
rect 183652 608398 183704 608404
rect 193692 608394 193720 610028
rect 204916 608394 204944 632062
rect 212368 629898 212396 632266
rect 221372 632256 221424 632262
rect 221372 632198 221424 632204
rect 212060 629870 212396 629898
rect 221384 629898 221412 632198
rect 232596 632188 232648 632194
rect 232596 632130 232648 632136
rect 231032 632120 231084 632126
rect 231032 632062 231084 632068
rect 232504 632120 232556 632126
rect 232504 632062 232556 632068
rect 231044 629898 231072 632062
rect 221384 629870 221720 629898
rect 231044 629870 231380 629898
rect 209686 620256 209742 620265
rect 209686 620191 209742 620200
rect 205638 619576 205694 619585
rect 205638 619511 205694 619520
rect 205652 611250 205680 619511
rect 209700 611318 209728 620191
rect 209688 611312 209740 611318
rect 209688 611254 209740 611260
rect 205640 611244 205692 611250
rect 205640 611186 205692 611192
rect 231676 611244 231728 611250
rect 231676 611186 231728 611192
rect 231688 610722 231716 611186
rect 231380 610694 231716 610722
rect 211724 610014 212060 610042
rect 221720 610014 222056 610042
rect 211724 608462 211752 610014
rect 222028 608462 222056 610014
rect 232516 608462 232544 632062
rect 232608 611250 232636 632130
rect 232700 611998 232728 632266
rect 233238 619576 233294 619585
rect 233238 619511 233294 619520
rect 232688 611992 232740 611998
rect 232688 611934 232740 611940
rect 232596 611244 232648 611250
rect 232596 611186 232648 611192
rect 233252 611182 233280 619511
rect 233240 611176 233292 611182
rect 233240 611118 233292 611124
rect 211712 608456 211764 608462
rect 211712 608398 211764 608404
rect 222016 608456 222068 608462
rect 222016 608398 222068 608404
rect 232504 608456 232556 608462
rect 232504 608398 232556 608404
rect 81992 608388 82044 608394
rect 81992 608330 82044 608336
rect 95884 608388 95936 608394
rect 95884 608330 95936 608336
rect 99472 608388 99524 608394
rect 99472 608330 99524 608336
rect 109684 608388 109736 608394
rect 109684 608330 109736 608336
rect 120724 608388 120776 608394
rect 120724 608330 120776 608336
rect 127072 608388 127124 608394
rect 127072 608330 127124 608336
rect 137652 608388 137704 608394
rect 137652 608330 137704 608336
rect 148416 608388 148468 608394
rect 148416 608330 148468 608336
rect 193680 608388 193732 608394
rect 193680 608330 193732 608336
rect 204904 608388 204956 608394
rect 204904 608330 204956 608336
rect 119436 604716 119488 604722
rect 119436 604658 119488 604664
rect 137652 604716 137704 604722
rect 137652 604658 137704 604664
rect 148324 604716 148376 604722
rect 148324 604658 148376 604664
rect 165712 604716 165764 604722
rect 165712 604658 165764 604664
rect 175464 604716 175516 604722
rect 175464 604658 175516 604664
rect 193680 604716 193732 604722
rect 193680 604658 193732 604664
rect 203524 604716 203576 604722
rect 203524 604658 203576 604664
rect 221372 604716 221424 604722
rect 221372 604658 221424 604664
rect 81440 604648 81492 604654
rect 81440 604590 81492 604596
rect 91468 604648 91520 604654
rect 91468 604590 91520 604596
rect 109684 604648 109736 604654
rect 109684 604590 109736 604596
rect 81452 602970 81480 604590
rect 91100 604580 91152 604586
rect 91100 604522 91152 604528
rect 91112 602970 91140 604522
rect 81452 602942 81696 602970
rect 91112 602942 91356 602970
rect 71884 602262 72036 602290
rect 71044 580916 71096 580922
rect 71044 580858 71096 580864
rect 71884 580854 71912 602262
rect 91480 583794 91508 604590
rect 94504 604580 94556 604586
rect 94504 604522 94556 604528
rect 93858 592648 93914 592657
rect 93858 592583 93914 592592
rect 91356 583766 91508 583794
rect 93872 583642 93900 592583
rect 93860 583636 93912 583642
rect 93860 583578 93912 583584
rect 72036 583086 72096 583114
rect 81696 583086 82032 583114
rect 71872 580848 71924 580854
rect 71872 580790 71924 580796
rect 72068 580786 72096 583086
rect 82004 580786 82032 583086
rect 94516 580786 94544 604522
rect 109696 602956 109724 604590
rect 119344 604580 119396 604586
rect 119344 604522 119396 604528
rect 119356 602956 119384 604522
rect 99484 602262 100050 602290
rect 97906 593328 97962 593337
rect 97906 593263 97962 593272
rect 97920 583642 97948 593263
rect 97908 583636 97960 583642
rect 97908 583578 97960 583584
rect 99484 580786 99512 602262
rect 119448 583794 119476 604658
rect 127992 604648 128044 604654
rect 127992 604590 128044 604596
rect 120724 604580 120776 604586
rect 120724 604522 120776 604528
rect 119370 583766 119476 583794
rect 100036 580854 100064 583100
rect 100024 580848 100076 580854
rect 100024 580790 100076 580796
rect 109696 580786 109724 583100
rect 120736 580786 120764 604522
rect 128004 602956 128032 604590
rect 137664 602956 137692 604658
rect 147312 604580 147364 604586
rect 147312 604522 147364 604528
rect 147324 602956 147352 604522
rect 126886 593328 126942 593337
rect 126886 593263 126942 593272
rect 121458 592648 121514 592657
rect 121458 592583 121514 592592
rect 121472 583710 121500 592583
rect 126900 583710 126928 593263
rect 148336 586514 148364 604658
rect 148508 604648 148560 604654
rect 148508 604590 148560 604596
rect 156328 604648 156380 604654
rect 156328 604590 156380 604596
rect 148416 604580 148468 604586
rect 148416 604522 148468 604528
rect 147784 586486 148364 586514
rect 121460 583704 121512 583710
rect 121460 583646 121512 583652
rect 126888 583704 126940 583710
rect 147784 583658 147812 586486
rect 126888 583646 126940 583652
rect 147338 583630 147812 583658
rect 128004 580854 128032 583100
rect 137664 580854 137692 583100
rect 148428 580854 148456 604522
rect 148520 584458 148548 604590
rect 156340 602970 156368 604590
rect 156032 602942 156368 602970
rect 165724 602834 165752 604658
rect 175372 604580 175424 604586
rect 175372 604522 175424 604528
rect 175384 602834 175412 604522
rect 165692 602806 165752 602834
rect 175352 602806 175412 602834
rect 154486 593328 154542 593337
rect 154486 593263 154542 593272
rect 149058 592648 149114 592657
rect 149058 592583 149114 592592
rect 148508 584452 148560 584458
rect 148508 584394 148560 584400
rect 149072 583642 149100 592583
rect 154500 583642 154528 593263
rect 155868 584452 155920 584458
rect 155868 584394 155920 584400
rect 155880 583794 155908 584394
rect 175476 583794 175504 604658
rect 178684 604648 178736 604654
rect 178684 604590 178736 604596
rect 177304 604580 177356 604586
rect 177304 604522 177356 604528
rect 155880 583766 156032 583794
rect 175352 583766 175504 583794
rect 149060 583636 149112 583642
rect 149060 583578 149112 583584
rect 154488 583636 154540 583642
rect 154488 583578 154540 583584
rect 165692 583086 166028 583114
rect 166000 580854 166028 583086
rect 177316 580854 177344 604522
rect 178038 592648 178094 592657
rect 178038 592583 178094 592592
rect 178052 583710 178080 592583
rect 178040 583704 178092 583710
rect 178040 583646 178092 583652
rect 178696 580990 178724 604590
rect 193692 602956 193720 604658
rect 203340 604580 203392 604586
rect 203340 604522 203392 604528
rect 203352 602956 203380 604522
rect 183664 602262 184046 602290
rect 182086 593328 182142 593337
rect 182086 593263 182142 593272
rect 182100 583574 182128 593263
rect 182088 583568 182140 583574
rect 182088 583510 182140 583516
rect 178684 580984 178736 580990
rect 178684 580926 178736 580932
rect 183664 580854 183692 602262
rect 203536 583794 203564 604658
rect 204904 604580 204956 604586
rect 204904 604522 204956 604528
rect 203366 583766 203564 583794
rect 184032 580990 184060 583100
rect 184020 580984 184072 580990
rect 184020 580926 184072 580932
rect 127992 580848 128044 580854
rect 127992 580790 128044 580796
rect 137652 580848 137704 580854
rect 137652 580790 137704 580796
rect 148416 580848 148468 580854
rect 148416 580790 148468 580796
rect 165988 580848 166040 580854
rect 165988 580790 166040 580796
rect 177304 580848 177356 580854
rect 177304 580790 177356 580796
rect 183652 580848 183704 580854
rect 183652 580790 183704 580796
rect 193692 580786 193720 583100
rect 204916 580786 204944 604522
rect 212356 604512 212408 604518
rect 212356 604454 212408 604460
rect 212368 602970 212396 604454
rect 212060 602942 212396 602970
rect 221384 602970 221412 604658
rect 232504 604648 232556 604654
rect 232504 604590 232556 604596
rect 231032 604580 231084 604586
rect 231032 604522 231084 604528
rect 231044 602970 231072 604522
rect 221384 602942 221720 602970
rect 231044 602942 231380 602970
rect 209686 593328 209742 593337
rect 209686 593263 209742 593272
rect 205638 592648 205694 592657
rect 205638 592583 205694 592592
rect 205652 583642 205680 592583
rect 209700 583710 209728 593263
rect 232516 586514 232544 604590
rect 232596 604580 232648 604586
rect 232596 604522 232648 604528
rect 231872 586486 232544 586514
rect 209688 583704 209740 583710
rect 231872 583658 231900 586486
rect 209688 583646 209740 583652
rect 205640 583636 205692 583642
rect 231380 583630 231900 583658
rect 205640 583578 205692 583584
rect 211724 583086 212060 583114
rect 221720 583086 222056 583114
rect 211724 580854 211752 583086
rect 222028 580854 222056 583086
rect 232608 580854 232636 604522
rect 232688 604512 232740 604518
rect 232688 604454 232740 604460
rect 232700 584458 232728 604454
rect 233238 592648 233294 592657
rect 233238 592583 233294 592592
rect 232688 584452 232740 584458
rect 232688 584394 232740 584400
rect 233252 583574 233280 592583
rect 233240 583568 233292 583574
rect 233240 583510 233292 583516
rect 211712 580848 211764 580854
rect 211712 580790 211764 580796
rect 222016 580848 222068 580854
rect 222016 580790 222068 580796
rect 232596 580848 232648 580854
rect 232596 580790 232648 580796
rect 72056 580780 72108 580786
rect 72056 580722 72108 580728
rect 81992 580780 82044 580786
rect 81992 580722 82044 580728
rect 94504 580780 94556 580786
rect 94504 580722 94556 580728
rect 99472 580780 99524 580786
rect 99472 580722 99524 580728
rect 109684 580780 109736 580786
rect 109684 580722 109736 580728
rect 120724 580780 120776 580786
rect 120724 580722 120776 580728
rect 193680 580780 193732 580786
rect 193680 580722 193732 580728
rect 204904 580780 204956 580786
rect 204904 580722 204956 580728
rect 71044 578468 71096 578474
rect 71044 578410 71096 578416
rect 69664 578264 69716 578270
rect 69664 578206 69716 578212
rect 69676 554606 69704 578206
rect 70306 566264 70362 566273
rect 70306 566199 70362 566208
rect 70320 557394 70348 566199
rect 70308 557388 70360 557394
rect 70308 557330 70360 557336
rect 69664 554600 69716 554606
rect 69664 554542 69716 554548
rect 70306 539336 70362 539345
rect 70306 539271 70362 539280
rect 70320 529786 70348 539271
rect 70308 529780 70360 529786
rect 70308 529722 70360 529728
rect 71056 527066 71084 578410
rect 148416 578400 148468 578406
rect 148416 578342 148468 578348
rect 165620 578400 165672 578406
rect 165620 578342 165672 578348
rect 175464 578400 175516 578406
rect 175464 578342 175516 578348
rect 193680 578400 193732 578406
rect 193680 578342 193732 578348
rect 203524 578400 203576 578406
rect 203524 578342 203576 578348
rect 221372 578400 221424 578406
rect 221372 578342 221424 578348
rect 232504 578400 232556 578406
rect 232504 578342 232556 578348
rect 81440 578332 81492 578338
rect 81440 578274 81492 578280
rect 91468 578332 91520 578338
rect 91468 578274 91520 578280
rect 109684 578332 109736 578338
rect 109684 578274 109736 578280
rect 119436 578332 119488 578338
rect 119436 578274 119488 578280
rect 137652 578332 137704 578338
rect 137652 578274 137704 578280
rect 81452 575906 81480 578274
rect 91100 578264 91152 578270
rect 91100 578206 91152 578212
rect 91112 575906 91140 578206
rect 81452 575878 81696 575906
rect 91112 575878 91356 575906
rect 71884 575334 72036 575362
rect 71884 554674 71912 575334
rect 91480 556730 91508 578274
rect 94504 578264 94556 578270
rect 94504 578206 94556 578212
rect 93858 565584 93914 565593
rect 93858 565519 93914 565528
rect 93872 557462 93900 565519
rect 93860 557456 93912 557462
rect 93860 557398 93912 557404
rect 91356 556702 91508 556730
rect 72036 556022 72096 556050
rect 81696 556022 82032 556050
rect 72068 554742 72096 556022
rect 72056 554736 72108 554742
rect 72056 554678 72108 554684
rect 71872 554668 71924 554674
rect 71872 554610 71924 554616
rect 82004 554606 82032 556022
rect 94516 554606 94544 578206
rect 109696 575892 109724 578274
rect 119344 578264 119396 578270
rect 119344 578206 119396 578212
rect 119356 575892 119384 578206
rect 99484 575334 100050 575362
rect 97906 566264 97962 566273
rect 97906 566199 97962 566208
rect 97920 557530 97948 566199
rect 97908 557524 97960 557530
rect 97908 557466 97960 557472
rect 99484 554742 99512 575334
rect 119448 556730 119476 578274
rect 120724 578264 120776 578270
rect 120724 578206 120776 578212
rect 119370 556702 119476 556730
rect 99472 554736 99524 554742
rect 99472 554678 99524 554684
rect 100036 554674 100064 556036
rect 100024 554668 100076 554674
rect 100024 554610 100076 554616
rect 109696 554606 109724 556036
rect 120736 554606 120764 578206
rect 137664 575892 137692 578274
rect 147312 578264 147364 578270
rect 147312 578206 147364 578212
rect 148324 578264 148376 578270
rect 148324 578206 148376 578212
rect 147324 575892 147352 578206
rect 127084 575334 128018 575362
rect 126886 566264 126942 566273
rect 126886 566199 126942 566208
rect 121458 565584 121514 565593
rect 121458 565519 121514 565528
rect 121472 557394 121500 565519
rect 126900 557462 126928 566199
rect 126888 557456 126940 557462
rect 126888 557398 126940 557404
rect 121460 557388 121512 557394
rect 121460 557330 121512 557336
rect 127084 554742 127112 575334
rect 147680 562352 147732 562358
rect 147680 562294 147732 562300
rect 147692 556730 147720 562294
rect 147338 556702 147720 556730
rect 127072 554736 127124 554742
rect 127072 554678 127124 554684
rect 128004 554674 128032 556036
rect 127992 554668 128044 554674
rect 127992 554610 128044 554616
rect 137664 554606 137692 556036
rect 148336 554606 148364 578206
rect 148428 562358 148456 578342
rect 156328 578332 156380 578338
rect 156328 578274 156380 578280
rect 156340 575906 156368 578274
rect 165632 576178 165660 578342
rect 175280 578264 175332 578270
rect 175280 578206 175332 578212
rect 175292 576178 175320 578206
rect 165632 576150 165706 576178
rect 175292 576150 175366 576178
rect 156032 575878 156368 575906
rect 165678 575892 165706 576150
rect 175338 575892 175366 576150
rect 154486 566264 154542 566273
rect 154486 566199 154542 566208
rect 149058 565584 149114 565593
rect 149058 565519 149114 565528
rect 148416 562352 148468 562358
rect 148416 562294 148468 562300
rect 149072 557530 149100 565519
rect 154500 557530 154528 566199
rect 149060 557524 149112 557530
rect 149060 557466 149112 557472
rect 154488 557524 154540 557530
rect 154488 557466 154540 557472
rect 175476 556730 175504 578342
rect 178684 578332 178736 578338
rect 178684 578274 178736 578280
rect 177304 578264 177356 578270
rect 177304 578206 177356 578212
rect 175352 556702 175504 556730
rect 156032 556022 156092 556050
rect 165692 556022 166028 556050
rect 156064 554674 156092 556022
rect 166000 554674 166028 556022
rect 177316 554674 177344 578206
rect 178038 565584 178094 565593
rect 178038 565519 178094 565528
rect 178052 557462 178080 565519
rect 178040 557456 178092 557462
rect 178040 557398 178092 557404
rect 178696 554674 178724 578274
rect 193692 575892 193720 578342
rect 203340 578264 203392 578270
rect 203340 578206 203392 578212
rect 203352 575892 203380 578206
rect 183664 575334 184046 575362
rect 182086 566264 182142 566273
rect 182086 566199 182142 566208
rect 182100 557462 182128 566199
rect 182088 557456 182140 557462
rect 182088 557398 182140 557404
rect 183664 554742 183692 575334
rect 203536 556730 203564 578342
rect 212264 578332 212316 578338
rect 212264 578274 212316 578280
rect 204904 578264 204956 578270
rect 204904 578206 204956 578212
rect 203366 556702 203564 556730
rect 183652 554736 183704 554742
rect 183652 554678 183704 554684
rect 184032 554674 184060 556036
rect 156052 554668 156104 554674
rect 156052 554610 156104 554616
rect 165988 554668 166040 554674
rect 165988 554610 166040 554616
rect 177304 554668 177356 554674
rect 177304 554610 177356 554616
rect 178684 554668 178736 554674
rect 178684 554610 178736 554616
rect 184020 554668 184072 554674
rect 184020 554610 184072 554616
rect 193692 554606 193720 556036
rect 204916 554606 204944 578206
rect 212276 575906 212304 578274
rect 212060 575878 212304 575906
rect 221384 575906 221412 578342
rect 231032 578264 231084 578270
rect 231032 578206 231084 578212
rect 231044 575906 231072 578206
rect 221384 575878 221720 575906
rect 231044 575878 231380 575906
rect 209686 566264 209742 566273
rect 209686 566199 209742 566208
rect 205638 565584 205694 565593
rect 205638 565519 205694 565528
rect 205652 557530 205680 565519
rect 209700 557530 209728 566199
rect 232516 557534 232544 578342
rect 232688 578332 232740 578338
rect 232688 578274 232740 578280
rect 232596 578264 232648 578270
rect 232596 578206 232648 578212
rect 205640 557524 205692 557530
rect 205640 557466 205692 557472
rect 209688 557524 209740 557530
rect 209688 557466 209740 557472
rect 231780 557506 232544 557534
rect 231780 556730 231808 557506
rect 231380 556702 231808 556730
rect 211724 556022 212060 556050
rect 221720 556022 222056 556050
rect 211724 554674 211752 556022
rect 222028 554674 222056 556022
rect 232608 554674 232636 578206
rect 232700 558210 232728 578274
rect 233238 565584 233294 565593
rect 233238 565519 233294 565528
rect 232688 558204 232740 558210
rect 232688 558146 232740 558152
rect 233252 557462 233280 565519
rect 233240 557456 233292 557462
rect 233240 557398 233292 557404
rect 211712 554668 211764 554674
rect 211712 554610 211764 554616
rect 222016 554668 222068 554674
rect 222016 554610 222068 554616
rect 232596 554668 232648 554674
rect 232596 554610 232648 554616
rect 81992 554600 82044 554606
rect 81992 554542 82044 554548
rect 94504 554600 94556 554606
rect 94504 554542 94556 554548
rect 109684 554600 109736 554606
rect 109684 554542 109736 554548
rect 120724 554600 120776 554606
rect 120724 554542 120776 554548
rect 137652 554600 137704 554606
rect 137652 554542 137704 554548
rect 148324 554600 148376 554606
rect 148324 554542 148376 554548
rect 193680 554600 193732 554606
rect 193680 554542 193732 554548
rect 204904 554600 204956 554606
rect 204904 554542 204956 554548
rect 148324 550860 148376 550866
rect 148324 550802 148376 550808
rect 165712 550860 165764 550866
rect 165712 550802 165764 550808
rect 175464 550860 175516 550866
rect 175464 550802 175516 550808
rect 193680 550860 193732 550866
rect 193680 550802 193732 550808
rect 203524 550860 203576 550866
rect 203524 550802 203576 550808
rect 221372 550860 221424 550866
rect 221372 550802 221424 550808
rect 81440 550792 81492 550798
rect 81440 550734 81492 550740
rect 91468 550792 91520 550798
rect 91468 550734 91520 550740
rect 109684 550792 109736 550798
rect 109684 550734 109736 550740
rect 119436 550792 119488 550798
rect 119436 550734 119488 550740
rect 137652 550792 137704 550798
rect 137652 550734 137704 550740
rect 81452 548978 81480 550734
rect 91100 550724 91152 550730
rect 91100 550666 91152 550672
rect 91112 548978 91140 550666
rect 81452 548950 81696 548978
rect 91112 548950 91356 548978
rect 71884 548270 72036 548298
rect 71044 527060 71096 527066
rect 71044 527002 71096 527008
rect 71884 526998 71912 548270
rect 91480 529666 91508 550734
rect 94504 550724 94556 550730
rect 94504 550666 94556 550672
rect 93858 538656 93914 538665
rect 93858 538591 93914 538600
rect 93872 529854 93900 538591
rect 93860 529848 93912 529854
rect 93860 529790 93912 529796
rect 91356 529638 91508 529666
rect 72022 528850 72050 529108
rect 81696 529094 82032 529122
rect 71976 528822 72050 528850
rect 71872 526992 71924 526998
rect 71872 526934 71924 526940
rect 71976 526930 72004 528822
rect 82004 526930 82032 529094
rect 94516 526930 94544 550666
rect 109696 548964 109724 550734
rect 119344 550724 119396 550730
rect 119344 550666 119396 550672
rect 119356 548964 119384 550666
rect 99484 548270 100050 548298
rect 97906 539336 97962 539345
rect 97906 539271 97962 539280
rect 97920 529922 97948 539271
rect 97908 529916 97960 529922
rect 97908 529858 97960 529864
rect 99484 526930 99512 548270
rect 119448 529666 119476 550734
rect 120724 550724 120776 550730
rect 120724 550666 120776 550672
rect 119370 529638 119476 529666
rect 100036 526998 100064 529108
rect 100024 526992 100076 526998
rect 100024 526934 100076 526940
rect 109696 526930 109724 529108
rect 120736 526930 120764 550666
rect 137664 548964 137692 550734
rect 147312 550724 147364 550730
rect 147312 550666 147364 550672
rect 147324 548964 147352 550666
rect 127084 548270 128018 548298
rect 126886 539336 126942 539345
rect 126886 539271 126942 539280
rect 121458 538656 121514 538665
rect 121458 538591 121514 538600
rect 121472 529786 121500 538591
rect 126900 529854 126928 539271
rect 126888 529848 126940 529854
rect 126888 529790 126940 529796
rect 121460 529780 121512 529786
rect 121460 529722 121512 529728
rect 127084 526930 127112 548270
rect 148336 538214 148364 550802
rect 156328 550792 156380 550798
rect 156328 550734 156380 550740
rect 148416 550724 148468 550730
rect 148416 550666 148468 550672
rect 147784 538186 148364 538214
rect 147784 529666 147812 538186
rect 147338 529638 147812 529666
rect 128004 526998 128032 529108
rect 127992 526992 128044 526998
rect 127992 526934 128044 526940
rect 137664 526930 137692 529108
rect 148428 526930 148456 550666
rect 156340 548978 156368 550734
rect 156032 548950 156368 548978
rect 165724 548842 165752 550802
rect 175372 550724 175424 550730
rect 175372 550666 175424 550672
rect 175384 548842 175412 550666
rect 165692 548814 165752 548842
rect 175352 548814 175412 548842
rect 154486 539336 154542 539345
rect 154486 539271 154542 539280
rect 149058 538656 149114 538665
rect 149058 538591 149114 538600
rect 149072 529922 149100 538591
rect 154500 529922 154528 539271
rect 149060 529916 149112 529922
rect 149060 529858 149112 529864
rect 154488 529916 154540 529922
rect 154488 529858 154540 529864
rect 175476 529666 175504 550802
rect 178684 550792 178736 550798
rect 178684 550734 178736 550740
rect 177304 550724 177356 550730
rect 177304 550666 177356 550672
rect 175352 529638 175504 529666
rect 156018 528850 156046 529108
rect 165692 529094 166028 529122
rect 155972 528822 156046 528850
rect 155972 526998 156000 528822
rect 166000 526998 166028 529094
rect 177316 526998 177344 550666
rect 178038 538656 178094 538665
rect 178038 538591 178094 538600
rect 178052 529854 178080 538591
rect 178040 529848 178092 529854
rect 178040 529790 178092 529796
rect 178696 527134 178724 550734
rect 193692 548964 193720 550802
rect 203340 550724 203392 550730
rect 203340 550666 203392 550672
rect 203352 548964 203380 550666
rect 183664 548270 184046 548298
rect 182086 539336 182142 539345
rect 182086 539271 182142 539280
rect 182100 529854 182128 539271
rect 182088 529848 182140 529854
rect 182088 529790 182140 529796
rect 178684 527128 178736 527134
rect 178684 527070 178736 527076
rect 183664 526998 183692 548270
rect 203536 529666 203564 550802
rect 204904 550724 204956 550730
rect 204904 550666 204956 550672
rect 203366 529638 203564 529666
rect 184032 527134 184060 529108
rect 184020 527128 184072 527134
rect 184020 527070 184072 527076
rect 155960 526992 156012 526998
rect 155960 526934 156012 526940
rect 165988 526992 166040 526998
rect 165988 526934 166040 526940
rect 177304 526992 177356 526998
rect 177304 526934 177356 526940
rect 183652 526992 183704 526998
rect 183652 526934 183704 526940
rect 193692 526930 193720 529108
rect 204916 526930 204944 550666
rect 212356 550656 212408 550662
rect 212356 550598 212408 550604
rect 212368 548978 212396 550598
rect 212060 548950 212396 548978
rect 221384 548978 221412 550802
rect 232504 550792 232556 550798
rect 232504 550734 232556 550740
rect 231032 550724 231084 550730
rect 231032 550666 231084 550672
rect 231044 548978 231072 550666
rect 221384 548950 221720 548978
rect 231044 548950 231380 548978
rect 209686 539336 209742 539345
rect 209686 539271 209742 539280
rect 205638 538656 205694 538665
rect 205638 538591 205694 538600
rect 205652 529922 205680 538591
rect 209700 529922 209728 539271
rect 232516 538214 232544 550734
rect 232596 550724 232648 550730
rect 232596 550666 232648 550672
rect 231872 538186 232544 538214
rect 205640 529916 205692 529922
rect 205640 529858 205692 529864
rect 209688 529916 209740 529922
rect 209688 529858 209740 529864
rect 231872 529802 231900 538186
rect 231780 529774 231900 529802
rect 231780 529666 231808 529774
rect 231380 529638 231808 529666
rect 211724 529094 212060 529122
rect 221720 529094 221964 529122
rect 211724 526998 211752 529094
rect 221936 526998 221964 529094
rect 232608 526998 232636 550666
rect 232688 550656 232740 550662
rect 232688 550598 232740 550604
rect 232700 530262 232728 550598
rect 233238 538656 233294 538665
rect 233238 538591 233294 538600
rect 232688 530256 232740 530262
rect 232688 530198 232740 530204
rect 233252 529854 233280 538591
rect 233240 529848 233292 529854
rect 233240 529790 233292 529796
rect 211712 526992 211764 526998
rect 211712 526934 211764 526940
rect 221924 526992 221976 526998
rect 221924 526934 221976 526940
rect 232596 526992 232648 526998
rect 232596 526934 232648 526940
rect 71964 526924 72016 526930
rect 71964 526866 72016 526872
rect 81992 526924 82044 526930
rect 81992 526866 82044 526872
rect 94504 526924 94556 526930
rect 94504 526866 94556 526872
rect 99472 526924 99524 526930
rect 99472 526866 99524 526872
rect 109684 526924 109736 526930
rect 109684 526866 109736 526872
rect 120724 526924 120776 526930
rect 120724 526866 120776 526872
rect 127072 526924 127124 526930
rect 127072 526866 127124 526872
rect 137652 526924 137704 526930
rect 137652 526866 137704 526872
rect 148416 526924 148468 526930
rect 148416 526866 148468 526872
rect 193680 526924 193732 526930
rect 193680 526866 193732 526872
rect 204904 526924 204956 526930
rect 204904 526866 204956 526872
rect 71044 523252 71096 523258
rect 71044 523194 71096 523200
rect 212356 523252 212408 523258
rect 212356 523194 212408 523200
rect 232688 523252 232740 523258
rect 232688 523194 232740 523200
rect 69664 523048 69716 523054
rect 69664 522990 69716 522996
rect 69676 500818 69704 522990
rect 70308 520328 70360 520334
rect 70308 520270 70360 520276
rect 70320 512281 70348 520270
rect 70306 512272 70362 512281
rect 70306 512207 70362 512216
rect 69664 500812 69716 500818
rect 69664 500754 69716 500760
rect 70306 484800 70362 484809
rect 70306 484735 70362 484744
rect 70320 476066 70348 484735
rect 70308 476060 70360 476066
rect 70308 476002 70360 476008
rect 71056 473278 71084 523194
rect 148416 523184 148468 523190
rect 148416 523126 148468 523132
rect 165712 523184 165764 523190
rect 165712 523126 165764 523132
rect 175464 523184 175516 523190
rect 175464 523126 175516 523132
rect 193680 523184 193732 523190
rect 193680 523126 193732 523132
rect 203524 523184 203576 523190
rect 203524 523126 203576 523132
rect 81440 523116 81492 523122
rect 81440 523058 81492 523064
rect 91468 523116 91520 523122
rect 91468 523058 91520 523064
rect 109684 523116 109736 523122
rect 109684 523058 109736 523064
rect 119436 523116 119488 523122
rect 119436 523058 119488 523064
rect 137652 523116 137704 523122
rect 137652 523058 137704 523064
rect 81452 521914 81480 523058
rect 91100 523048 91152 523054
rect 91100 522990 91152 522996
rect 91112 521914 91140 522990
rect 81452 521886 81696 521914
rect 91112 521886 91356 521914
rect 71884 521206 72036 521234
rect 71884 500886 71912 521206
rect 91480 502738 91508 523058
rect 94504 523048 94556 523054
rect 94504 522990 94556 522996
rect 93860 520396 93912 520402
rect 93860 520338 93912 520344
rect 93872 511601 93900 520338
rect 93858 511592 93914 511601
rect 93858 511527 93914 511536
rect 91356 502710 91508 502738
rect 72036 502030 72096 502058
rect 81696 502030 82032 502058
rect 72068 500954 72096 502030
rect 72056 500948 72108 500954
rect 72056 500890 72108 500896
rect 71872 500880 71924 500886
rect 71872 500822 71924 500828
rect 82004 500818 82032 502030
rect 94516 500818 94544 522990
rect 109696 521900 109724 523058
rect 119344 523048 119396 523054
rect 119344 522990 119396 522996
rect 119356 521900 119384 522990
rect 99484 521206 100050 521234
rect 97906 512272 97962 512281
rect 97906 512207 97962 512216
rect 97920 503674 97948 512207
rect 97908 503668 97960 503674
rect 97908 503610 97960 503616
rect 99484 500954 99512 521206
rect 119448 502738 119476 523058
rect 120724 523048 120776 523054
rect 120724 522990 120776 522996
rect 119370 502710 119476 502738
rect 99472 500948 99524 500954
rect 99472 500890 99524 500896
rect 100036 500886 100064 502044
rect 100024 500880 100076 500886
rect 100024 500822 100076 500828
rect 109696 500818 109724 502044
rect 120736 500818 120764 522990
rect 137664 521900 137692 523058
rect 147312 523048 147364 523054
rect 147312 522990 147364 522996
rect 148324 523048 148376 523054
rect 148324 522990 148376 522996
rect 147324 521900 147352 522990
rect 127084 521206 128018 521234
rect 121460 520328 121512 520334
rect 121460 520270 121512 520276
rect 126888 520328 126940 520334
rect 126888 520270 126940 520276
rect 121472 511601 121500 520270
rect 126900 512281 126928 520270
rect 126886 512272 126942 512281
rect 126886 512207 126942 512216
rect 121458 511592 121514 511601
rect 121458 511527 121514 511536
rect 127084 500954 127112 521206
rect 147680 505640 147732 505646
rect 147680 505582 147732 505588
rect 147692 502738 147720 505582
rect 147338 502710 147720 502738
rect 127072 500948 127124 500954
rect 127072 500890 127124 500896
rect 128004 500886 128032 502044
rect 127992 500880 128044 500886
rect 127992 500822 128044 500828
rect 137664 500818 137692 502044
rect 148336 500818 148364 522990
rect 148428 505646 148456 523126
rect 156328 523116 156380 523122
rect 156328 523058 156380 523064
rect 156340 521914 156368 523058
rect 156032 521886 156368 521914
rect 165724 521778 165752 523126
rect 175372 523048 175424 523054
rect 175372 522990 175424 522996
rect 175384 521778 175412 522990
rect 165692 521750 165752 521778
rect 175352 521750 175412 521778
rect 155868 520396 155920 520402
rect 155868 520338 155920 520344
rect 155880 518906 155908 520338
rect 154488 518900 154540 518906
rect 154488 518842 154540 518848
rect 155868 518900 155920 518906
rect 155868 518842 155920 518848
rect 154500 512281 154528 518842
rect 154486 512272 154542 512281
rect 154486 512207 154542 512216
rect 149058 511592 149114 511601
rect 149058 511527 149114 511536
rect 148416 505640 148468 505646
rect 148416 505582 148468 505588
rect 149072 503674 149100 511527
rect 149060 503668 149112 503674
rect 149060 503610 149112 503616
rect 175476 502738 175504 523126
rect 178684 523116 178736 523122
rect 178684 523058 178736 523064
rect 177304 523048 177356 523054
rect 177304 522990 177356 522996
rect 175352 502710 175504 502738
rect 156032 502030 156092 502058
rect 165692 502030 166028 502058
rect 156064 500886 156092 502030
rect 166000 500886 166028 502030
rect 177316 500886 177344 522990
rect 178040 520328 178092 520334
rect 178040 520270 178092 520276
rect 178052 511601 178080 520270
rect 178038 511592 178094 511601
rect 178038 511527 178094 511536
rect 178696 500886 178724 523058
rect 193692 521900 193720 523126
rect 203340 523048 203392 523054
rect 203340 522990 203392 522996
rect 203352 521900 203380 522990
rect 183664 521206 184046 521234
rect 182086 512272 182142 512281
rect 182086 512207 182142 512216
rect 182100 503674 182128 512207
rect 182088 503668 182140 503674
rect 182088 503610 182140 503616
rect 183664 500954 183692 521206
rect 203536 502738 203564 523126
rect 204904 523048 204956 523054
rect 204904 522990 204956 522996
rect 203366 502710 203564 502738
rect 183652 500948 183704 500954
rect 183652 500890 183704 500896
rect 184032 500886 184060 502044
rect 156052 500880 156104 500886
rect 156052 500822 156104 500828
rect 165988 500880 166040 500886
rect 165988 500822 166040 500828
rect 177304 500880 177356 500886
rect 177304 500822 177356 500828
rect 178684 500880 178736 500886
rect 178684 500822 178736 500828
rect 184020 500880 184072 500886
rect 184020 500822 184072 500828
rect 193692 500818 193720 502044
rect 204916 500818 204944 522990
rect 212368 521914 212396 523194
rect 221372 523184 221424 523190
rect 221372 523126 221424 523132
rect 212060 521886 212396 521914
rect 221384 521914 221412 523126
rect 232504 523116 232556 523122
rect 232504 523058 232556 523064
rect 231032 523048 231084 523054
rect 231032 522990 231084 522996
rect 231044 521914 231072 522990
rect 221384 521886 221720 521914
rect 231044 521886 231380 521914
rect 205640 520396 205692 520402
rect 205640 520338 205692 520344
rect 205652 511601 205680 520338
rect 209688 520328 209740 520334
rect 209688 520270 209740 520276
rect 209700 512281 209728 520270
rect 209686 512272 209742 512281
rect 209686 512207 209742 512216
rect 205638 511592 205694 511601
rect 205638 511527 205694 511536
rect 232516 509234 232544 523058
rect 232596 523048 232648 523054
rect 232596 522990 232648 522996
rect 231872 509206 232544 509234
rect 231872 502874 231900 509206
rect 231780 502846 231900 502874
rect 231780 502738 231808 502846
rect 231380 502710 231808 502738
rect 211724 502030 212060 502058
rect 221720 502030 222056 502058
rect 211724 500886 211752 502030
rect 222028 500886 222056 502030
rect 232608 500886 232636 522990
rect 232700 504286 232728 523194
rect 233238 511592 233294 511601
rect 233238 511527 233294 511536
rect 232688 504280 232740 504286
rect 232688 504222 232740 504228
rect 233252 503674 233280 511527
rect 233240 503668 233292 503674
rect 233240 503610 233292 503616
rect 211712 500880 211764 500886
rect 211712 500822 211764 500828
rect 222016 500880 222068 500886
rect 222016 500822 222068 500828
rect 232596 500880 232648 500886
rect 232596 500822 232648 500828
rect 81992 500812 82044 500818
rect 81992 500754 82044 500760
rect 94504 500812 94556 500818
rect 94504 500754 94556 500760
rect 109684 500812 109736 500818
rect 109684 500754 109736 500760
rect 120724 500812 120776 500818
rect 120724 500754 120776 500760
rect 137652 500812 137704 500818
rect 137652 500754 137704 500760
rect 148324 500812 148376 500818
rect 148324 500754 148376 500760
rect 193680 500812 193732 500818
rect 193680 500754 193732 500760
rect 204904 500812 204956 500818
rect 204904 500754 204956 500760
rect 148416 497072 148468 497078
rect 148416 497014 148468 497020
rect 165712 497072 165764 497078
rect 165712 497014 165764 497020
rect 175464 497072 175516 497078
rect 175464 497014 175516 497020
rect 193680 497072 193732 497078
rect 193680 497014 193732 497020
rect 203524 497072 203576 497078
rect 203524 497014 203576 497020
rect 221372 497072 221424 497078
rect 221372 497014 221424 497020
rect 81440 497004 81492 497010
rect 81440 496946 81492 496952
rect 91468 497004 91520 497010
rect 91468 496946 91520 496952
rect 109684 497004 109736 497010
rect 109684 496946 109736 496952
rect 119436 497004 119488 497010
rect 119436 496946 119488 496952
rect 137652 497004 137704 497010
rect 137652 496946 137704 496952
rect 81452 494986 81480 496946
rect 91100 496936 91152 496942
rect 91100 496878 91152 496884
rect 91112 494986 91140 496878
rect 81452 494958 81696 494986
rect 91112 494958 91356 494986
rect 71884 494278 72036 494306
rect 71044 473272 71096 473278
rect 71044 473214 71096 473220
rect 71884 473210 71912 494278
rect 91480 475674 91508 496946
rect 94504 496936 94556 496942
rect 94504 496878 94556 496884
rect 93858 484664 93914 484673
rect 93858 484599 93914 484608
rect 93872 475998 93900 484599
rect 93860 475992 93912 475998
rect 93860 475934 93912 475940
rect 91356 475646 91508 475674
rect 72036 475102 72096 475130
rect 81696 475102 82032 475130
rect 71872 473204 71924 473210
rect 71872 473146 71924 473152
rect 72068 473142 72096 475102
rect 82004 473142 82032 475102
rect 94516 473142 94544 496878
rect 109696 494972 109724 496946
rect 119344 496936 119396 496942
rect 119344 496878 119396 496884
rect 119356 494972 119384 496878
rect 99484 494278 100050 494306
rect 97906 485344 97962 485353
rect 97906 485279 97962 485288
rect 97920 475998 97948 485279
rect 97908 475992 97960 475998
rect 97908 475934 97960 475940
rect 99484 473142 99512 494278
rect 119448 475674 119476 496946
rect 120724 496936 120776 496942
rect 120724 496878 120776 496884
rect 119370 475646 119476 475674
rect 100036 473210 100064 475116
rect 100024 473204 100076 473210
rect 100024 473146 100076 473152
rect 109696 473142 109724 475116
rect 120736 473142 120764 496878
rect 137664 494972 137692 496946
rect 147312 496936 147364 496942
rect 147312 496878 147364 496884
rect 148324 496936 148376 496942
rect 148324 496878 148376 496884
rect 147324 494972 147352 496878
rect 127084 494278 128018 494306
rect 126886 485344 126942 485353
rect 126886 485279 126942 485288
rect 121458 484664 121514 484673
rect 121458 484599 121514 484608
rect 121472 476066 121500 484599
rect 126900 476066 126928 485279
rect 121460 476060 121512 476066
rect 121460 476002 121512 476008
rect 126888 476060 126940 476066
rect 126888 476002 126940 476008
rect 127084 473142 127112 494278
rect 147680 477692 147732 477698
rect 147680 477634 147732 477640
rect 147692 475674 147720 477634
rect 147338 475646 147720 475674
rect 128004 473210 128032 475116
rect 127992 473204 128044 473210
rect 127992 473146 128044 473152
rect 137664 473142 137692 475116
rect 148336 473142 148364 496878
rect 148428 477698 148456 497014
rect 156328 497004 156380 497010
rect 156328 496946 156380 496952
rect 156340 494986 156368 496946
rect 156032 494958 156368 494986
rect 165724 494850 165752 497014
rect 175372 496936 175424 496942
rect 175372 496878 175424 496884
rect 175384 494850 175412 496878
rect 165692 494822 165752 494850
rect 175352 494822 175412 494850
rect 154486 485344 154542 485353
rect 154486 485279 154542 485288
rect 149058 484664 149114 484673
rect 149058 484599 149114 484608
rect 148416 477692 148468 477698
rect 148416 477634 148468 477640
rect 149072 475998 149100 484599
rect 154500 475998 154528 485279
rect 149060 475992 149112 475998
rect 149060 475934 149112 475940
rect 154488 475992 154540 475998
rect 154488 475934 154540 475940
rect 175476 475674 175504 497014
rect 178684 497004 178736 497010
rect 178684 496946 178736 496952
rect 177304 496936 177356 496942
rect 177304 496878 177356 496884
rect 175352 475646 175504 475674
rect 156032 475102 156092 475130
rect 165692 475102 166028 475130
rect 156064 473210 156092 475102
rect 166000 473210 166028 475102
rect 177316 473210 177344 496878
rect 178038 484664 178094 484673
rect 178038 484599 178094 484608
rect 178052 476066 178080 484599
rect 178040 476060 178092 476066
rect 178040 476002 178092 476008
rect 178696 473346 178724 496946
rect 193692 494972 193720 497014
rect 203340 496936 203392 496942
rect 203340 496878 203392 496884
rect 203352 494972 203380 496878
rect 183664 494278 184046 494306
rect 182086 485344 182142 485353
rect 182086 485279 182142 485288
rect 182100 475930 182128 485279
rect 182088 475924 182140 475930
rect 182088 475866 182140 475872
rect 178684 473340 178736 473346
rect 178684 473282 178736 473288
rect 183664 473210 183692 494278
rect 203536 475674 203564 497014
rect 204904 496936 204956 496942
rect 204904 496878 204956 496884
rect 203366 475646 203564 475674
rect 184032 473346 184060 475116
rect 184020 473340 184072 473346
rect 184020 473282 184072 473288
rect 156052 473204 156104 473210
rect 156052 473146 156104 473152
rect 165988 473204 166040 473210
rect 165988 473146 166040 473152
rect 177304 473204 177356 473210
rect 177304 473146 177356 473152
rect 183652 473204 183704 473210
rect 183652 473146 183704 473152
rect 193692 473142 193720 475116
rect 204916 473142 204944 496878
rect 212356 496868 212408 496874
rect 212356 496810 212408 496816
rect 212368 494986 212396 496810
rect 212060 494958 212396 494986
rect 221384 494986 221412 497014
rect 232504 497004 232556 497010
rect 232504 496946 232556 496952
rect 231032 496936 231084 496942
rect 231032 496878 231084 496884
rect 231044 494986 231072 496878
rect 221384 494958 221720 494986
rect 231044 494958 231380 494986
rect 209686 485344 209742 485353
rect 209686 485279 209742 485288
rect 205638 484528 205694 484537
rect 205638 484463 205694 484472
rect 205652 475998 205680 484463
rect 209700 476066 209728 485279
rect 232516 480254 232544 496946
rect 232596 496936 232648 496942
rect 232596 496878 232648 496884
rect 231872 480226 232544 480254
rect 209688 476060 209740 476066
rect 209688 476002 209740 476008
rect 205640 475992 205692 475998
rect 205640 475934 205692 475940
rect 231872 475810 231900 480226
rect 231780 475782 231900 475810
rect 231780 475674 231808 475782
rect 231380 475646 231808 475674
rect 211724 475102 212060 475130
rect 221720 475102 222056 475130
rect 211724 473210 211752 475102
rect 222028 473210 222056 475102
rect 232608 473210 232636 496878
rect 232688 496868 232740 496874
rect 232688 496810 232740 496816
rect 232700 476610 232728 496810
rect 233238 484664 233294 484673
rect 233238 484599 233294 484608
rect 232688 476604 232740 476610
rect 232688 476546 232740 476552
rect 233252 475930 233280 484599
rect 233240 475924 233292 475930
rect 233240 475866 233292 475872
rect 211712 473204 211764 473210
rect 211712 473146 211764 473152
rect 222016 473204 222068 473210
rect 222016 473146 222068 473152
rect 232596 473204 232648 473210
rect 232596 473146 232648 473152
rect 72056 473136 72108 473142
rect 72056 473078 72108 473084
rect 81992 473136 82044 473142
rect 81992 473078 82044 473084
rect 94504 473136 94556 473142
rect 94504 473078 94556 473084
rect 99472 473136 99524 473142
rect 99472 473078 99524 473084
rect 109684 473136 109736 473142
rect 109684 473078 109736 473084
rect 120724 473136 120776 473142
rect 120724 473078 120776 473084
rect 127072 473136 127124 473142
rect 127072 473078 127124 473084
rect 137652 473136 137704 473142
rect 137652 473078 137704 473084
rect 148324 473136 148376 473142
rect 148324 473078 148376 473084
rect 193680 473136 193732 473142
rect 193680 473078 193732 473084
rect 204904 473136 204956 473142
rect 204904 473078 204956 473084
rect 71044 469464 71096 469470
rect 71044 469406 71096 469412
rect 69664 469260 69716 469266
rect 69664 469202 69716 469208
rect 69676 445602 69704 469202
rect 70308 466472 70360 466478
rect 70308 466414 70360 466420
rect 70320 458289 70348 466414
rect 70306 458280 70362 458289
rect 70306 458215 70362 458224
rect 69664 445596 69716 445602
rect 69664 445538 69716 445544
rect 69664 443216 69716 443222
rect 69664 443158 69716 443164
rect 69676 391882 69704 443158
rect 70306 430808 70362 430817
rect 70306 430743 70362 430752
rect 70320 422278 70348 430743
rect 70308 422272 70360 422278
rect 70308 422214 70360 422220
rect 71056 419422 71084 469406
rect 148416 469396 148468 469402
rect 148416 469338 148468 469344
rect 165712 469396 165764 469402
rect 165712 469338 165764 469344
rect 175464 469396 175516 469402
rect 175464 469338 175516 469344
rect 193680 469396 193732 469402
rect 193680 469338 193732 469344
rect 203524 469396 203576 469402
rect 203524 469338 203576 469344
rect 221372 469396 221424 469402
rect 221372 469338 221424 469344
rect 232504 469396 232556 469402
rect 232504 469338 232556 469344
rect 81440 469328 81492 469334
rect 81440 469270 81492 469276
rect 91468 469328 91520 469334
rect 91468 469270 91520 469276
rect 109684 469328 109736 469334
rect 109684 469270 109736 469276
rect 119436 469328 119488 469334
rect 119436 469270 119488 469276
rect 137652 469328 137704 469334
rect 137652 469270 137704 469276
rect 81452 467922 81480 469270
rect 91100 469260 91152 469266
rect 91100 469202 91152 469208
rect 91112 467922 91140 469202
rect 81452 467894 81696 467922
rect 91112 467894 91356 467922
rect 71884 467214 72036 467242
rect 71884 445670 71912 467214
rect 91480 448746 91508 469270
rect 94504 469260 94556 469266
rect 94504 469202 94556 469208
rect 93860 466540 93912 466546
rect 93860 466482 93912 466488
rect 93872 457609 93900 466482
rect 93858 457600 93914 457609
rect 93858 457535 93914 457544
rect 91356 448718 91508 448746
rect 72036 448038 72096 448066
rect 81696 448038 82032 448066
rect 72068 445738 72096 448038
rect 72056 445732 72108 445738
rect 72056 445674 72108 445680
rect 71872 445664 71924 445670
rect 71872 445606 71924 445612
rect 82004 445602 82032 448038
rect 94516 445602 94544 469202
rect 109696 467908 109724 469270
rect 119344 469260 119396 469266
rect 119344 469202 119396 469208
rect 119356 467908 119384 469202
rect 99484 467214 100050 467242
rect 97908 466540 97960 466546
rect 97908 466482 97960 466488
rect 97920 458289 97948 466482
rect 97906 458280 97962 458289
rect 97906 458215 97962 458224
rect 99484 445738 99512 467214
rect 119448 448746 119476 469270
rect 120724 469260 120776 469266
rect 120724 469202 120776 469208
rect 119370 448718 119476 448746
rect 99472 445732 99524 445738
rect 99472 445674 99524 445680
rect 100036 445670 100064 448052
rect 100024 445664 100076 445670
rect 100024 445606 100076 445612
rect 109696 445602 109724 448052
rect 120736 445602 120764 469202
rect 137664 467908 137692 469270
rect 147312 469260 147364 469266
rect 147312 469202 147364 469208
rect 148324 469260 148376 469266
rect 148324 469202 148376 469208
rect 147324 467908 147352 469202
rect 127084 467214 128018 467242
rect 121460 466472 121512 466478
rect 121460 466414 121512 466420
rect 126888 466472 126940 466478
rect 126888 466414 126940 466420
rect 121472 457609 121500 466414
rect 126900 458289 126928 466414
rect 126886 458280 126942 458289
rect 126886 458215 126942 458224
rect 121458 457600 121514 457609
rect 121458 457535 121514 457544
rect 127084 445738 127112 467214
rect 147680 448520 147732 448526
rect 147338 448468 147680 448474
rect 147338 448462 147732 448468
rect 147338 448446 147720 448462
rect 127072 445732 127124 445738
rect 127072 445674 127124 445680
rect 128004 445670 128032 448052
rect 127992 445664 128044 445670
rect 127992 445606 128044 445612
rect 137664 445602 137692 448052
rect 148336 445602 148364 469202
rect 148428 448526 148456 469338
rect 156328 469328 156380 469334
rect 156328 469270 156380 469276
rect 156340 467922 156368 469270
rect 156032 467894 156368 467922
rect 165724 467786 165752 469338
rect 175372 469260 175424 469266
rect 175372 469202 175424 469208
rect 175384 467786 175412 469202
rect 165692 467758 165752 467786
rect 175352 467758 175412 467786
rect 149060 466540 149112 466546
rect 149060 466482 149112 466488
rect 154488 466540 154540 466546
rect 154488 466482 154540 466488
rect 149072 457609 149100 466482
rect 154500 458289 154528 466482
rect 154486 458280 154542 458289
rect 154486 458215 154542 458224
rect 149058 457600 149114 457609
rect 149058 457535 149114 457544
rect 175476 448746 175504 469338
rect 178684 469328 178736 469334
rect 178684 469270 178736 469276
rect 177304 469260 177356 469266
rect 177304 469202 177356 469208
rect 175352 448718 175504 448746
rect 148416 448520 148468 448526
rect 148416 448462 148468 448468
rect 156032 448038 156092 448066
rect 165692 448038 166028 448066
rect 156064 445670 156092 448038
rect 166000 445670 166028 448038
rect 177316 445670 177344 469202
rect 178040 466472 178092 466478
rect 178040 466414 178092 466420
rect 178052 457609 178080 466414
rect 178038 457600 178094 457609
rect 178038 457535 178094 457544
rect 178696 445670 178724 469270
rect 193692 467908 193720 469338
rect 203340 469260 203392 469266
rect 203340 469202 203392 469208
rect 203352 467908 203380 469202
rect 183664 467214 184046 467242
rect 182088 466608 182140 466614
rect 182088 466550 182140 466556
rect 182100 458289 182128 466550
rect 182086 458280 182142 458289
rect 182086 458215 182142 458224
rect 183664 445738 183692 467214
rect 203536 448746 203564 469338
rect 212356 469328 212408 469334
rect 212356 469270 212408 469276
rect 204904 469260 204956 469266
rect 204904 469202 204956 469208
rect 203366 448718 203564 448746
rect 183652 445732 183704 445738
rect 183652 445674 183704 445680
rect 184032 445670 184060 448052
rect 156052 445664 156104 445670
rect 156052 445606 156104 445612
rect 165988 445664 166040 445670
rect 165988 445606 166040 445612
rect 177304 445664 177356 445670
rect 177304 445606 177356 445612
rect 178684 445664 178736 445670
rect 178684 445606 178736 445612
rect 184020 445664 184072 445670
rect 184020 445606 184072 445612
rect 193692 445602 193720 448052
rect 204916 445602 204944 469202
rect 212368 467922 212396 469270
rect 212060 467894 212396 467922
rect 221384 467922 221412 469338
rect 231032 469260 231084 469266
rect 231032 469202 231084 469208
rect 231044 467922 231072 469202
rect 221384 467894 221720 467922
rect 231044 467894 231380 467922
rect 205640 466540 205692 466546
rect 205640 466482 205692 466488
rect 205652 457609 205680 466482
rect 209688 466472 209740 466478
rect 209688 466414 209740 466420
rect 209700 458289 209728 466414
rect 209686 458280 209742 458289
rect 209686 458215 209742 458224
rect 205638 457600 205694 457609
rect 205638 457535 205694 457544
rect 232516 451274 232544 469338
rect 232688 469328 232740 469334
rect 232688 469270 232740 469276
rect 232596 469260 232648 469266
rect 232596 469202 232648 469208
rect 231872 451246 232544 451274
rect 231872 448474 231900 451246
rect 231380 448446 231900 448474
rect 211724 448038 212060 448066
rect 221720 448038 222056 448066
rect 211724 445670 211752 448038
rect 222028 445670 222056 448038
rect 232608 445670 232636 469202
rect 232700 449954 232728 469270
rect 233240 466608 233292 466614
rect 233240 466550 233292 466556
rect 233252 457609 233280 466550
rect 233238 457600 233294 457609
rect 233238 457535 233294 457544
rect 232688 449948 232740 449954
rect 232688 449890 232740 449896
rect 211712 445664 211764 445670
rect 211712 445606 211764 445612
rect 222016 445664 222068 445670
rect 222016 445606 222068 445612
rect 232596 445664 232648 445670
rect 232596 445606 232648 445612
rect 81992 445596 82044 445602
rect 81992 445538 82044 445544
rect 94504 445596 94556 445602
rect 94504 445538 94556 445544
rect 109684 445596 109736 445602
rect 109684 445538 109736 445544
rect 120724 445596 120776 445602
rect 120724 445538 120776 445544
rect 137652 445596 137704 445602
rect 137652 445538 137704 445544
rect 148324 445596 148376 445602
rect 148324 445538 148376 445544
rect 193680 445596 193732 445602
rect 193680 445538 193732 445544
rect 204904 445596 204956 445602
rect 204904 445538 204956 445544
rect 212264 443216 212316 443222
rect 212264 443158 212316 443164
rect 232688 443216 232740 443222
rect 232688 443158 232740 443164
rect 81440 443148 81492 443154
rect 81440 443090 81492 443096
rect 148324 443148 148376 443154
rect 148324 443090 148376 443096
rect 165620 443148 165672 443154
rect 165620 443090 165672 443096
rect 175464 443148 175516 443154
rect 175464 443090 175516 443096
rect 193680 443148 193732 443154
rect 193680 443090 193732 443096
rect 203524 443148 203576 443154
rect 203524 443090 203576 443096
rect 81452 440994 81480 443090
rect 91100 443080 91152 443086
rect 91100 443022 91152 443028
rect 91468 443080 91520 443086
rect 91468 443022 91520 443028
rect 109684 443080 109736 443086
rect 109684 443022 109736 443028
rect 119436 443080 119488 443086
rect 119436 443022 119488 443028
rect 137284 443080 137336 443086
rect 137284 443022 137336 443028
rect 91112 440994 91140 443022
rect 81452 440966 81696 440994
rect 91112 440966 91356 440994
rect 71884 440286 72036 440314
rect 71044 419416 71096 419422
rect 71044 419358 71096 419364
rect 71884 419354 71912 440286
rect 91480 421682 91508 443022
rect 94504 443012 94556 443018
rect 94504 442954 94556 442960
rect 93860 440292 93912 440298
rect 93860 440234 93912 440240
rect 93872 430681 93900 440234
rect 93858 430672 93914 430681
rect 93858 430607 93914 430616
rect 91356 421654 91508 421682
rect 72036 421110 72096 421138
rect 81696 421110 82032 421138
rect 71872 419348 71924 419354
rect 71872 419290 71924 419296
rect 72068 419286 72096 421110
rect 82004 419286 82032 421110
rect 94516 419286 94544 442954
rect 109696 440980 109724 443022
rect 119344 443012 119396 443018
rect 119344 442954 119396 442960
rect 119356 440980 119384 442954
rect 97908 440292 97960 440298
rect 97908 440234 97960 440240
rect 99484 440286 100050 440314
rect 97920 431361 97948 440234
rect 97906 431352 97962 431361
rect 97906 431287 97962 431296
rect 99484 419286 99512 440286
rect 119448 421682 119476 443022
rect 120724 443012 120776 443018
rect 120724 442954 120776 442960
rect 119370 421654 119476 421682
rect 100036 419354 100064 421124
rect 100024 419348 100076 419354
rect 100024 419290 100076 419296
rect 109696 419286 109724 421124
rect 120736 419286 120764 442954
rect 137296 440994 137324 443022
rect 147036 443012 147088 443018
rect 147036 442954 147088 442960
rect 147048 440994 147076 442954
rect 137296 440966 137678 440994
rect 147048 440966 147338 440994
rect 127084 440286 128018 440314
rect 126886 431352 126942 431361
rect 126886 431287 126942 431296
rect 121458 430672 121514 430681
rect 121458 430607 121514 430616
rect 121472 422278 121500 430607
rect 126900 422278 126928 431287
rect 121460 422272 121512 422278
rect 121460 422214 121512 422220
rect 126888 422272 126940 422278
rect 126888 422214 126940 422220
rect 127084 419286 127112 440286
rect 148336 422294 148364 443090
rect 156328 443080 156380 443086
rect 156328 443022 156380 443028
rect 148416 443012 148468 443018
rect 148416 442954 148468 442960
rect 147784 422266 148364 422294
rect 147784 421682 147812 422266
rect 147338 421654 147812 421682
rect 128004 419354 128032 421124
rect 127992 419348 128044 419354
rect 127992 419290 128044 419296
rect 137664 419286 137692 421124
rect 148428 419286 148456 442954
rect 156340 440994 156368 443022
rect 165632 441130 165660 443090
rect 175280 443012 175332 443018
rect 175280 442954 175332 442960
rect 175292 441130 175320 442954
rect 165632 441102 165706 441130
rect 175292 441102 175366 441130
rect 156032 440966 156368 440994
rect 165678 440980 165706 441102
rect 175338 440980 175366 441102
rect 149060 440292 149112 440298
rect 149060 440234 149112 440240
rect 154488 440292 154540 440298
rect 154488 440234 154540 440240
rect 149072 430681 149100 440234
rect 154500 431361 154528 440234
rect 154486 431352 154542 431361
rect 154486 431287 154542 431296
rect 149058 430672 149114 430681
rect 149058 430607 149114 430616
rect 175476 421682 175504 443090
rect 178684 443080 178736 443086
rect 178684 443022 178736 443028
rect 177304 443012 177356 443018
rect 177304 442954 177356 442960
rect 175352 421654 175504 421682
rect 156032 421110 156092 421138
rect 165692 421110 166028 421138
rect 156064 419354 156092 421110
rect 166000 419354 166028 421110
rect 177316 419354 177344 442954
rect 178038 430672 178094 430681
rect 178038 430607 178094 430616
rect 178052 422278 178080 430607
rect 178040 422272 178092 422278
rect 178040 422214 178092 422220
rect 178696 419490 178724 443022
rect 193692 440980 193720 443090
rect 203340 443012 203392 443018
rect 203340 442954 203392 442960
rect 203352 440980 203380 442954
rect 182088 440360 182140 440366
rect 182088 440302 182140 440308
rect 182100 431361 182128 440302
rect 183664 440286 184046 440314
rect 182086 431352 182142 431361
rect 182086 431287 182142 431296
rect 178684 419484 178736 419490
rect 178684 419426 178736 419432
rect 183664 419354 183692 440286
rect 203536 421682 203564 443090
rect 204904 443012 204956 443018
rect 204904 442954 204956 442960
rect 203366 421654 203564 421682
rect 184032 419490 184060 421124
rect 184020 419484 184072 419490
rect 184020 419426 184072 419432
rect 156052 419348 156104 419354
rect 156052 419290 156104 419296
rect 165988 419348 166040 419354
rect 165988 419290 166040 419296
rect 177304 419348 177356 419354
rect 177304 419290 177356 419296
rect 183652 419348 183704 419354
rect 183652 419290 183704 419296
rect 193692 419286 193720 421124
rect 204916 419286 204944 442954
rect 212276 440994 212304 443158
rect 221372 443148 221424 443154
rect 221372 443090 221424 443096
rect 212060 440966 212304 440994
rect 221384 440994 221412 443090
rect 232504 443080 232556 443086
rect 232504 443022 232556 443028
rect 231032 443012 231084 443018
rect 231032 442954 231084 442960
rect 231044 440994 231072 442954
rect 221384 440966 221720 440994
rect 231044 440966 231380 440994
rect 205640 440292 205692 440298
rect 205640 440234 205692 440240
rect 205652 431225 205680 440234
rect 209686 431352 209742 431361
rect 209686 431287 209742 431296
rect 205638 431216 205694 431225
rect 205638 431151 205694 431160
rect 209700 422278 209728 431287
rect 232516 422294 232544 443022
rect 232596 443012 232648 443018
rect 232596 442954 232648 442960
rect 209688 422272 209740 422278
rect 209688 422214 209740 422220
rect 231780 422266 232544 422294
rect 231780 421682 231808 422266
rect 231380 421654 231808 421682
rect 211724 421110 212060 421138
rect 221720 421110 222056 421138
rect 211724 419354 211752 421110
rect 222028 419354 222056 421110
rect 232608 419354 232636 442954
rect 232700 423026 232728 443158
rect 233240 440360 233292 440366
rect 233240 440302 233292 440308
rect 233252 430681 233280 440302
rect 233238 430672 233294 430681
rect 233238 430607 233294 430616
rect 232688 423020 232740 423026
rect 232688 422962 232740 422968
rect 211712 419348 211764 419354
rect 211712 419290 211764 419296
rect 222016 419348 222068 419354
rect 222016 419290 222068 419296
rect 232596 419348 232648 419354
rect 232596 419290 232648 419296
rect 72056 419280 72108 419286
rect 72056 419222 72108 419228
rect 81992 419280 82044 419286
rect 81992 419222 82044 419228
rect 94504 419280 94556 419286
rect 94504 419222 94556 419228
rect 99472 419280 99524 419286
rect 99472 419222 99524 419228
rect 109684 419280 109736 419286
rect 109684 419222 109736 419228
rect 120724 419280 120776 419286
rect 120724 419222 120776 419228
rect 127072 419280 127124 419286
rect 127072 419222 127124 419228
rect 137652 419280 137704 419286
rect 137652 419222 137704 419228
rect 148416 419280 148468 419286
rect 148416 419222 148468 419228
rect 193680 419280 193732 419286
rect 193680 419222 193732 419228
rect 204904 419280 204956 419286
rect 204904 419222 204956 419228
rect 119436 415676 119488 415682
rect 119436 415618 119488 415624
rect 137652 415676 137704 415682
rect 137652 415618 137704 415624
rect 148324 415676 148376 415682
rect 148324 415618 148376 415624
rect 165712 415676 165764 415682
rect 165712 415618 165764 415624
rect 175464 415676 175516 415682
rect 175464 415618 175516 415624
rect 193680 415676 193732 415682
rect 193680 415618 193732 415624
rect 203524 415676 203576 415682
rect 203524 415618 203576 415624
rect 221372 415676 221424 415682
rect 221372 415618 221424 415624
rect 81440 415608 81492 415614
rect 81440 415550 81492 415556
rect 91468 415608 91520 415614
rect 91468 415550 91520 415556
rect 109684 415608 109736 415614
rect 109684 415550 109736 415556
rect 81452 413930 81480 415550
rect 91100 415540 91152 415546
rect 91100 415482 91152 415488
rect 91112 413930 91140 415482
rect 81452 413902 81696 413930
rect 91112 413902 91356 413930
rect 71884 413222 72036 413250
rect 70306 404288 70362 404297
rect 70306 404223 70362 404232
rect 70320 394670 70348 404223
rect 70308 394664 70360 394670
rect 70308 394606 70360 394612
rect 69664 391876 69716 391882
rect 69664 391818 69716 391824
rect 71884 391814 71912 413222
rect 91480 394754 91508 415550
rect 94504 415540 94556 415546
rect 94504 415482 94556 415488
rect 93858 403608 93914 403617
rect 93858 403543 93914 403552
rect 91356 394726 91508 394754
rect 93872 394602 93900 403543
rect 93860 394596 93912 394602
rect 93860 394538 93912 394544
rect 72022 393802 72050 394060
rect 81696 394046 82032 394074
rect 71976 393774 72050 393802
rect 71872 391808 71924 391814
rect 71872 391750 71924 391756
rect 71976 391746 72004 393774
rect 82004 391746 82032 394046
rect 94516 391746 94544 415482
rect 109696 413916 109724 415550
rect 119344 415540 119396 415546
rect 119344 415482 119396 415488
rect 119356 413916 119384 415482
rect 99484 413222 100050 413250
rect 97906 404288 97962 404297
rect 97906 404223 97962 404232
rect 97920 394602 97948 404223
rect 97908 394596 97960 394602
rect 97908 394538 97960 394544
rect 99484 391746 99512 413222
rect 119448 394754 119476 415618
rect 127992 415608 128044 415614
rect 127992 415550 128044 415556
rect 120724 415540 120776 415546
rect 120724 415482 120776 415488
rect 119370 394726 119476 394754
rect 100036 391814 100064 394060
rect 100024 391808 100076 391814
rect 100024 391750 100076 391756
rect 109696 391746 109724 394060
rect 120736 391746 120764 415482
rect 128004 413916 128032 415550
rect 137664 413916 137692 415618
rect 147312 415540 147364 415546
rect 147312 415482 147364 415488
rect 147324 413916 147352 415482
rect 126886 404288 126942 404297
rect 126886 404223 126942 404232
rect 121458 403608 121514 403617
rect 121458 403543 121514 403552
rect 121472 394670 121500 403543
rect 126900 394670 126928 404223
rect 148336 402974 148364 415618
rect 148508 415608 148560 415614
rect 148508 415550 148560 415556
rect 156328 415608 156380 415614
rect 156328 415550 156380 415556
rect 148416 415540 148468 415546
rect 148416 415482 148468 415488
rect 147784 402946 148364 402974
rect 121460 394664 121512 394670
rect 121460 394606 121512 394612
rect 126888 394664 126940 394670
rect 147784 394618 147812 402946
rect 126888 394606 126940 394612
rect 147338 394590 147812 394618
rect 128004 391814 128032 394060
rect 137664 391814 137692 394060
rect 148428 391814 148456 415482
rect 148520 395350 148548 415550
rect 156340 413930 156368 415550
rect 156032 413902 156368 413930
rect 165724 413794 165752 415618
rect 175372 415540 175424 415546
rect 175372 415482 175424 415488
rect 175384 413794 175412 415482
rect 165692 413766 165752 413794
rect 175352 413766 175412 413794
rect 154486 404288 154542 404297
rect 154486 404223 154542 404232
rect 149058 403608 149114 403617
rect 149058 403543 149114 403552
rect 148508 395344 148560 395350
rect 148508 395286 148560 395292
rect 149072 394602 149100 403543
rect 149060 394596 149112 394602
rect 149060 394538 149112 394544
rect 154500 394534 154528 404223
rect 155868 395344 155920 395350
rect 155868 395286 155920 395292
rect 155880 394754 155908 395286
rect 175476 394754 175504 415618
rect 178684 415608 178736 415614
rect 178684 415550 178736 415556
rect 177304 415540 177356 415546
rect 177304 415482 177356 415488
rect 155880 394726 156032 394754
rect 175352 394726 175504 394754
rect 154488 394528 154540 394534
rect 154488 394470 154540 394476
rect 165692 394046 166028 394074
rect 166000 391814 166028 394046
rect 177316 391814 177344 415482
rect 178038 403608 178094 403617
rect 178038 403543 178094 403552
rect 178052 394670 178080 403543
rect 178040 394664 178092 394670
rect 178040 394606 178092 394612
rect 178696 391950 178724 415550
rect 193692 413916 193720 415618
rect 203340 415540 203392 415546
rect 203340 415482 203392 415488
rect 203352 413916 203380 415482
rect 183664 413222 184046 413250
rect 182086 404288 182142 404297
rect 182086 404223 182142 404232
rect 182100 394602 182128 404223
rect 182088 394596 182140 394602
rect 182088 394538 182140 394544
rect 178684 391944 178736 391950
rect 178684 391886 178736 391892
rect 183664 391814 183692 413222
rect 203536 394754 203564 415618
rect 204904 415540 204956 415546
rect 204904 415482 204956 415488
rect 203366 394726 203564 394754
rect 184032 391950 184060 394060
rect 184020 391944 184072 391950
rect 184020 391886 184072 391892
rect 127992 391808 128044 391814
rect 127992 391750 128044 391756
rect 137652 391808 137704 391814
rect 137652 391750 137704 391756
rect 148416 391808 148468 391814
rect 148416 391750 148468 391756
rect 165988 391808 166040 391814
rect 165988 391750 166040 391756
rect 177304 391808 177356 391814
rect 177304 391750 177356 391756
rect 183652 391808 183704 391814
rect 183652 391750 183704 391756
rect 193692 391746 193720 394060
rect 204916 391746 204944 415482
rect 212356 415472 212408 415478
rect 212356 415414 212408 415420
rect 212368 413930 212396 415414
rect 212060 413902 212396 413930
rect 221384 413930 221412 415618
rect 232596 415608 232648 415614
rect 232596 415550 232648 415556
rect 231032 415540 231084 415546
rect 231032 415482 231084 415488
rect 232504 415540 232556 415546
rect 232504 415482 232556 415488
rect 231044 413930 231072 415482
rect 221384 413902 221720 413930
rect 231044 413902 231380 413930
rect 209686 404288 209742 404297
rect 209686 404223 209742 404232
rect 205638 403608 205694 403617
rect 205638 403543 205694 403552
rect 205652 394534 205680 403543
rect 209700 394670 209728 404223
rect 209688 394664 209740 394670
rect 209688 394606 209740 394612
rect 205640 394528 205692 394534
rect 205640 394470 205692 394476
rect 211724 394046 212060 394074
rect 221720 394046 221964 394074
rect 231380 394046 231624 394074
rect 211724 391814 211752 394046
rect 221936 391814 221964 394046
rect 231596 393310 231624 394046
rect 231584 393304 231636 393310
rect 231584 393246 231636 393252
rect 232516 391814 232544 415482
rect 232608 393310 232636 415550
rect 232688 415472 232740 415478
rect 232688 415414 232740 415420
rect 232700 395078 232728 415414
rect 233238 403608 233294 403617
rect 233238 403543 233294 403552
rect 232688 395072 232740 395078
rect 232688 395014 232740 395020
rect 233252 394602 233280 403543
rect 233240 394596 233292 394602
rect 233240 394538 233292 394544
rect 232596 393304 232648 393310
rect 232596 393246 232648 393252
rect 211712 391808 211764 391814
rect 211712 391750 211764 391756
rect 221924 391808 221976 391814
rect 221924 391750 221976 391756
rect 232504 391808 232556 391814
rect 232504 391750 232556 391756
rect 71964 391740 72016 391746
rect 71964 391682 72016 391688
rect 81992 391740 82044 391746
rect 81992 391682 82044 391688
rect 94504 391740 94556 391746
rect 94504 391682 94556 391688
rect 99472 391740 99524 391746
rect 99472 391682 99524 391688
rect 109684 391740 109736 391746
rect 109684 391682 109736 391688
rect 120724 391740 120776 391746
rect 120724 391682 120776 391688
rect 193680 391740 193732 391746
rect 193680 391682 193732 391688
rect 204904 391740 204956 391746
rect 204904 391682 204956 391688
rect 71044 389428 71096 389434
rect 71044 389370 71096 389376
rect 212356 389428 212408 389434
rect 212356 389370 212408 389376
rect 232688 389428 232740 389434
rect 232688 389370 232740 389376
rect 69664 389224 69716 389230
rect 69664 389166 69716 389172
rect 69676 365566 69704 389166
rect 70306 376816 70362 376825
rect 70306 376751 70362 376760
rect 70320 368490 70348 376751
rect 70308 368484 70360 368490
rect 70308 368426 70360 368432
rect 69664 365560 69716 365566
rect 69664 365502 69716 365508
rect 70306 350296 70362 350305
rect 70306 350231 70362 350240
rect 70320 340882 70348 350231
rect 70308 340876 70360 340882
rect 70308 340818 70360 340824
rect 71056 338026 71084 389370
rect 148416 389360 148468 389366
rect 148416 389302 148468 389308
rect 165712 389360 165764 389366
rect 165712 389302 165764 389308
rect 175464 389360 175516 389366
rect 175464 389302 175516 389308
rect 193680 389360 193732 389366
rect 193680 389302 193732 389308
rect 203524 389360 203576 389366
rect 203524 389302 203576 389308
rect 81440 389292 81492 389298
rect 81440 389234 81492 389240
rect 91468 389292 91520 389298
rect 91468 389234 91520 389240
rect 109684 389292 109736 389298
rect 109684 389234 109736 389240
rect 119436 389292 119488 389298
rect 119436 389234 119488 389240
rect 137652 389292 137704 389298
rect 137652 389234 137704 389240
rect 81452 386866 81480 389234
rect 91100 389224 91152 389230
rect 91100 389166 91152 389172
rect 91112 386866 91140 389166
rect 81452 386838 81696 386866
rect 91112 386838 91356 386866
rect 71884 386294 72036 386322
rect 71884 365634 71912 386294
rect 91480 367690 91508 389234
rect 94504 389224 94556 389230
rect 94504 389166 94556 389172
rect 93858 376000 93914 376009
rect 93858 375935 93914 375944
rect 93872 368422 93900 375935
rect 93860 368416 93912 368422
rect 93860 368358 93912 368364
rect 91356 367662 91508 367690
rect 72036 367118 72096 367146
rect 81696 367118 82032 367146
rect 72068 365702 72096 367118
rect 72056 365696 72108 365702
rect 72056 365638 72108 365644
rect 71872 365628 71924 365634
rect 71872 365570 71924 365576
rect 82004 365566 82032 367118
rect 94516 365566 94544 389166
rect 109696 386852 109724 389234
rect 119344 389224 119396 389230
rect 119344 389166 119396 389172
rect 119356 386852 119384 389166
rect 99668 386294 100050 386322
rect 97906 376816 97962 376825
rect 97906 376751 97962 376760
rect 97920 368422 97948 376751
rect 99668 373994 99696 386294
rect 99484 373966 99696 373994
rect 97908 368416 97960 368422
rect 97908 368358 97960 368364
rect 99484 365702 99512 373966
rect 119448 367690 119476 389234
rect 120724 389224 120776 389230
rect 120724 389166 120776 389172
rect 119370 367662 119476 367690
rect 99472 365696 99524 365702
rect 99472 365638 99524 365644
rect 100036 365634 100064 367132
rect 100024 365628 100076 365634
rect 100024 365570 100076 365576
rect 109696 365566 109724 367132
rect 120736 365566 120764 389166
rect 137664 386852 137692 389234
rect 147312 389224 147364 389230
rect 147312 389166 147364 389172
rect 148324 389224 148376 389230
rect 148324 389166 148376 389172
rect 147324 386852 147352 389166
rect 127636 386294 128018 386322
rect 126886 376816 126942 376825
rect 126886 376751 126942 376760
rect 121458 376000 121514 376009
rect 121458 375935 121514 375944
rect 121472 368490 121500 375935
rect 126900 368490 126928 376751
rect 127636 373994 127664 386294
rect 127084 373966 127664 373994
rect 121460 368484 121512 368490
rect 121460 368426 121512 368432
rect 126888 368484 126940 368490
rect 126888 368426 126940 368432
rect 127084 365702 127112 373966
rect 147680 370592 147732 370598
rect 147680 370534 147732 370540
rect 147692 367690 147720 370534
rect 147338 367662 147720 367690
rect 127072 365696 127124 365702
rect 127072 365638 127124 365644
rect 128004 365634 128032 367132
rect 127992 365628 128044 365634
rect 127992 365570 128044 365576
rect 137664 365566 137692 367132
rect 148336 365566 148364 389166
rect 148428 370598 148456 389302
rect 156328 389292 156380 389298
rect 156328 389234 156380 389240
rect 156340 386866 156368 389234
rect 156032 386838 156368 386866
rect 165724 386730 165752 389302
rect 175372 389224 175424 389230
rect 175372 389166 175424 389172
rect 175384 386730 175412 389166
rect 165692 386702 165752 386730
rect 175352 386702 175412 386730
rect 154486 376816 154542 376825
rect 154486 376751 154542 376760
rect 149058 376000 149114 376009
rect 149058 375935 149114 375944
rect 148416 370592 148468 370598
rect 148416 370534 148468 370540
rect 149072 368422 149100 375935
rect 149060 368416 149112 368422
rect 149060 368358 149112 368364
rect 154500 368354 154528 376751
rect 154488 368348 154540 368354
rect 154488 368290 154540 368296
rect 175476 367690 175504 389302
rect 178684 389292 178736 389298
rect 178684 389234 178736 389240
rect 177304 389224 177356 389230
rect 177304 389166 177356 389172
rect 175352 367662 175504 367690
rect 156032 367118 156092 367146
rect 165692 367118 166028 367146
rect 156064 365634 156092 367118
rect 166000 365634 166028 367118
rect 177316 365634 177344 389166
rect 178038 376000 178094 376009
rect 178038 375935 178094 375944
rect 178052 368490 178080 375935
rect 178040 368484 178092 368490
rect 178040 368426 178092 368432
rect 178696 365634 178724 389234
rect 193692 386852 193720 389302
rect 203340 389224 203392 389230
rect 203340 389166 203392 389172
rect 203352 386852 203380 389166
rect 183664 386294 184046 386322
rect 182086 376816 182142 376825
rect 182086 376751 182142 376760
rect 182100 368422 182128 376751
rect 182088 368416 182140 368422
rect 182088 368358 182140 368364
rect 183664 365702 183692 386294
rect 203536 367690 203564 389302
rect 204904 389224 204956 389230
rect 204904 389166 204956 389172
rect 203366 367662 203564 367690
rect 183652 365696 183704 365702
rect 183652 365638 183704 365644
rect 184032 365634 184060 367132
rect 156052 365628 156104 365634
rect 156052 365570 156104 365576
rect 165988 365628 166040 365634
rect 165988 365570 166040 365576
rect 177304 365628 177356 365634
rect 177304 365570 177356 365576
rect 178684 365628 178736 365634
rect 178684 365570 178736 365576
rect 184020 365628 184072 365634
rect 184020 365570 184072 365576
rect 193692 365566 193720 367132
rect 204916 365566 204944 389166
rect 212368 386866 212396 389370
rect 221372 389360 221424 389366
rect 221372 389302 221424 389308
rect 212060 386838 212396 386866
rect 221384 386866 221412 389302
rect 232596 389292 232648 389298
rect 232596 389234 232648 389240
rect 231032 389224 231084 389230
rect 231032 389166 231084 389172
rect 232504 389224 232556 389230
rect 232504 389166 232556 389172
rect 231044 386866 231072 389166
rect 221384 386838 221720 386866
rect 231044 386838 231380 386866
rect 209686 377088 209742 377097
rect 209686 377023 209742 377032
rect 205638 376000 205694 376009
rect 205638 375935 205694 375944
rect 205652 368354 205680 375935
rect 209700 368490 209728 377023
rect 209688 368484 209740 368490
rect 209688 368426 209740 368432
rect 205640 368348 205692 368354
rect 205640 368290 205692 368296
rect 231676 368348 231728 368354
rect 231676 368290 231728 368296
rect 231688 367690 231716 368290
rect 231380 367662 231716 367690
rect 211724 367118 212060 367146
rect 221720 367118 222056 367146
rect 211724 365634 211752 367118
rect 222028 365634 222056 367118
rect 232516 365634 232544 389166
rect 232608 368354 232636 389234
rect 232700 369306 232728 389370
rect 233238 376000 233294 376009
rect 233238 375935 233294 375944
rect 232688 369300 232740 369306
rect 232688 369242 232740 369248
rect 233252 368422 233280 375935
rect 233240 368416 233292 368422
rect 233240 368358 233292 368364
rect 232596 368348 232648 368354
rect 232596 368290 232648 368296
rect 211712 365628 211764 365634
rect 211712 365570 211764 365576
rect 222016 365628 222068 365634
rect 222016 365570 222068 365576
rect 232504 365628 232556 365634
rect 232504 365570 232556 365576
rect 81992 365560 82044 365566
rect 81992 365502 82044 365508
rect 94504 365560 94556 365566
rect 94504 365502 94556 365508
rect 109684 365560 109736 365566
rect 109684 365502 109736 365508
rect 120724 365560 120776 365566
rect 120724 365502 120776 365508
rect 137652 365560 137704 365566
rect 137652 365502 137704 365508
rect 148324 365560 148376 365566
rect 148324 365502 148376 365508
rect 193680 365560 193732 365566
rect 193680 365502 193732 365508
rect 204904 365560 204956 365566
rect 204904 365502 204956 365508
rect 148416 361820 148468 361826
rect 148416 361762 148468 361768
rect 165712 361820 165764 361826
rect 165712 361762 165764 361768
rect 175464 361820 175516 361826
rect 175464 361762 175516 361768
rect 193680 361820 193732 361826
rect 193680 361762 193732 361768
rect 203524 361820 203576 361826
rect 203524 361762 203576 361768
rect 221372 361820 221424 361826
rect 221372 361762 221424 361768
rect 81440 361752 81492 361758
rect 81440 361694 81492 361700
rect 91468 361752 91520 361758
rect 91468 361694 91520 361700
rect 109684 361752 109736 361758
rect 109684 361694 109736 361700
rect 119436 361752 119488 361758
rect 119436 361694 119488 361700
rect 137652 361752 137704 361758
rect 137652 361694 137704 361700
rect 81452 359938 81480 361694
rect 91100 361684 91152 361690
rect 91100 361626 91152 361632
rect 91112 359938 91140 361626
rect 81452 359910 81696 359938
rect 91112 359910 91356 359938
rect 71884 359230 72036 359258
rect 71044 338020 71096 338026
rect 71044 337962 71096 337968
rect 71884 337958 71912 359230
rect 91480 340762 91508 361694
rect 94504 361684 94556 361690
rect 94504 361626 94556 361632
rect 93858 349616 93914 349625
rect 93858 349551 93914 349560
rect 93872 340814 93900 349551
rect 91356 340734 91508 340762
rect 93860 340808 93912 340814
rect 93860 340750 93912 340756
rect 72036 340054 72096 340082
rect 81696 340054 82032 340082
rect 71872 337952 71924 337958
rect 71872 337894 71924 337900
rect 72068 337890 72096 340054
rect 82004 337890 82032 340054
rect 94516 337890 94544 361626
rect 109696 359924 109724 361694
rect 119344 361684 119396 361690
rect 119344 361626 119396 361632
rect 119356 359924 119384 361626
rect 99484 359230 100050 359258
rect 97906 350296 97962 350305
rect 97906 350231 97962 350240
rect 97920 340814 97948 350231
rect 97908 340808 97960 340814
rect 97908 340750 97960 340756
rect 99484 337890 99512 359230
rect 119448 340762 119476 361694
rect 120724 361684 120776 361690
rect 120724 361626 120776 361632
rect 119370 340734 119476 340762
rect 100036 337958 100064 340068
rect 100024 337952 100076 337958
rect 100024 337894 100076 337900
rect 109696 337890 109724 340068
rect 120736 337890 120764 361626
rect 137664 359924 137692 361694
rect 147312 361684 147364 361690
rect 147312 361626 147364 361632
rect 148324 361684 148376 361690
rect 148324 361626 148376 361632
rect 147324 359924 147352 361626
rect 127084 359230 128018 359258
rect 126886 350296 126942 350305
rect 126886 350231 126942 350240
rect 121458 349616 121514 349625
rect 121458 349551 121514 349560
rect 121472 340882 121500 349551
rect 126900 340882 126928 350231
rect 121460 340876 121512 340882
rect 121460 340818 121512 340824
rect 126888 340876 126940 340882
rect 126888 340818 126940 340824
rect 127084 337890 127112 359230
rect 147680 342576 147732 342582
rect 147680 342518 147732 342524
rect 147692 340762 147720 342518
rect 147338 340734 147720 340762
rect 128004 337958 128032 340068
rect 127992 337952 128044 337958
rect 127992 337894 128044 337900
rect 137664 337890 137692 340068
rect 148336 337890 148364 361626
rect 148428 342582 148456 361762
rect 156328 361752 156380 361758
rect 156328 361694 156380 361700
rect 156340 359938 156368 361694
rect 156032 359910 156368 359938
rect 165724 359802 165752 361762
rect 175372 361684 175424 361690
rect 175372 361626 175424 361632
rect 175384 359802 175412 361626
rect 165692 359774 165752 359802
rect 175352 359774 175412 359802
rect 154486 350296 154542 350305
rect 154486 350231 154542 350240
rect 149058 349616 149114 349625
rect 149058 349551 149114 349560
rect 148416 342576 148468 342582
rect 148416 342518 148468 342524
rect 149072 340814 149100 349551
rect 154500 340814 154528 350231
rect 149060 340808 149112 340814
rect 149060 340750 149112 340756
rect 154488 340808 154540 340814
rect 175476 340762 175504 361762
rect 178684 361752 178736 361758
rect 178684 361694 178736 361700
rect 177304 361684 177356 361690
rect 177304 361626 177356 361632
rect 154488 340750 154540 340756
rect 175352 340734 175504 340762
rect 156032 340054 156092 340082
rect 165692 340054 166028 340082
rect 156064 337958 156092 340054
rect 166000 337958 166028 340054
rect 177316 337958 177344 361626
rect 178038 349616 178094 349625
rect 178038 349551 178094 349560
rect 178052 340882 178080 349551
rect 178040 340876 178092 340882
rect 178040 340818 178092 340824
rect 178696 338094 178724 361694
rect 193692 359924 193720 361762
rect 203340 361684 203392 361690
rect 203340 361626 203392 361632
rect 203352 359924 203380 361626
rect 183664 359230 184046 359258
rect 182086 350296 182142 350305
rect 182086 350231 182142 350240
rect 182100 340746 182128 350231
rect 182088 340740 182140 340746
rect 182088 340682 182140 340688
rect 178684 338088 178736 338094
rect 178684 338030 178736 338036
rect 183664 337958 183692 359230
rect 203536 340762 203564 361762
rect 204904 361684 204956 361690
rect 204904 361626 204956 361632
rect 203366 340734 203564 340762
rect 184032 338094 184060 340068
rect 184020 338088 184072 338094
rect 184020 338030 184072 338036
rect 156052 337952 156104 337958
rect 156052 337894 156104 337900
rect 165988 337952 166040 337958
rect 165988 337894 166040 337900
rect 177304 337952 177356 337958
rect 177304 337894 177356 337900
rect 183652 337952 183704 337958
rect 183652 337894 183704 337900
rect 193692 337890 193720 340068
rect 204916 337890 204944 361626
rect 212356 361616 212408 361622
rect 212356 361558 212408 361564
rect 212368 359938 212396 361558
rect 212060 359910 212396 359938
rect 221384 359938 221412 361762
rect 232596 361752 232648 361758
rect 232596 361694 232648 361700
rect 231032 361684 231084 361690
rect 231032 361626 231084 361632
rect 232504 361684 232556 361690
rect 232504 361626 232556 361632
rect 231044 359938 231072 361626
rect 221384 359910 221720 359938
rect 231044 359910 231380 359938
rect 209686 350296 209742 350305
rect 209686 350231 209742 350240
rect 205638 349616 205694 349625
rect 205638 349551 205694 349560
rect 205652 340814 205680 349551
rect 209700 340882 209728 350231
rect 209688 340876 209740 340882
rect 209688 340818 209740 340824
rect 205640 340808 205692 340814
rect 231676 340808 231728 340814
rect 205640 340750 205692 340756
rect 231380 340756 231676 340762
rect 231380 340750 231728 340756
rect 231380 340734 231716 340750
rect 211724 340054 212060 340082
rect 221720 340054 222056 340082
rect 211724 337958 211752 340054
rect 222028 337958 222056 340054
rect 232516 337958 232544 361626
rect 232608 340814 232636 361694
rect 232688 361616 232740 361622
rect 232688 361558 232740 361564
rect 232700 341426 232728 361558
rect 233238 349616 233294 349625
rect 233238 349551 233294 349560
rect 232688 341420 232740 341426
rect 232688 341362 232740 341368
rect 232596 340808 232648 340814
rect 232596 340750 232648 340756
rect 233252 340746 233280 349551
rect 233240 340740 233292 340746
rect 233240 340682 233292 340688
rect 211712 337952 211764 337958
rect 211712 337894 211764 337900
rect 222016 337952 222068 337958
rect 222016 337894 222068 337900
rect 232504 337952 232556 337958
rect 232504 337894 232556 337900
rect 72056 337884 72108 337890
rect 72056 337826 72108 337832
rect 81992 337884 82044 337890
rect 81992 337826 82044 337832
rect 94504 337884 94556 337890
rect 94504 337826 94556 337832
rect 99472 337884 99524 337890
rect 99472 337826 99524 337832
rect 109684 337884 109736 337890
rect 109684 337826 109736 337832
rect 120724 337884 120776 337890
rect 120724 337826 120776 337832
rect 127072 337884 127124 337890
rect 127072 337826 127124 337832
rect 137652 337884 137704 337890
rect 137652 337826 137704 337832
rect 148324 337884 148376 337890
rect 148324 337826 148376 337832
rect 193680 337884 193732 337890
rect 193680 337826 193732 337832
rect 204904 337884 204956 337890
rect 204904 337826 204956 337832
rect 71044 335572 71096 335578
rect 71044 335514 71096 335520
rect 212264 335572 212316 335578
rect 212264 335514 212316 335520
rect 232688 335572 232740 335578
rect 232688 335514 232740 335520
rect 69664 335368 69716 335374
rect 69664 335310 69716 335316
rect 69676 311710 69704 335310
rect 70306 322960 70362 322969
rect 70306 322895 70362 322904
rect 70320 314634 70348 322895
rect 70308 314628 70360 314634
rect 70308 314570 70360 314576
rect 69664 311704 69716 311710
rect 69664 311646 69716 311652
rect 70306 296304 70362 296313
rect 70306 296239 70362 296248
rect 70320 287026 70348 296239
rect 70308 287020 70360 287026
rect 70308 286962 70360 286968
rect 71056 284238 71084 335514
rect 148324 335504 148376 335510
rect 148324 335446 148376 335452
rect 165620 335504 165672 335510
rect 165620 335446 165672 335452
rect 175464 335504 175516 335510
rect 175464 335446 175516 335452
rect 193680 335504 193732 335510
rect 193680 335446 193732 335452
rect 203524 335504 203576 335510
rect 203524 335446 203576 335452
rect 81440 335436 81492 335442
rect 81440 335378 81492 335384
rect 91468 335436 91520 335442
rect 91468 335378 91520 335384
rect 109684 335436 109736 335442
rect 109684 335378 109736 335384
rect 119436 335436 119488 335442
rect 119436 335378 119488 335384
rect 137652 335436 137704 335442
rect 137652 335378 137704 335384
rect 81452 332874 81480 335378
rect 91100 335368 91152 335374
rect 91100 335310 91152 335316
rect 91112 332874 91140 335310
rect 81452 332846 81696 332874
rect 91112 332846 91356 332874
rect 71884 332302 72036 332330
rect 71884 311778 71912 332302
rect 91480 313698 91508 335378
rect 94504 335368 94556 335374
rect 94504 335310 94556 335316
rect 93858 322008 93914 322017
rect 93858 321943 93914 321952
rect 93872 314566 93900 321943
rect 93860 314560 93912 314566
rect 93860 314502 93912 314508
rect 91356 313670 91508 313698
rect 72036 313126 72096 313154
rect 81696 313126 82032 313154
rect 72068 311846 72096 313126
rect 72056 311840 72108 311846
rect 72056 311782 72108 311788
rect 71872 311772 71924 311778
rect 71872 311714 71924 311720
rect 82004 311710 82032 313126
rect 94516 311710 94544 335310
rect 109696 332860 109724 335378
rect 119344 335368 119396 335374
rect 119344 335310 119396 335316
rect 119356 332860 119384 335310
rect 99484 332302 100050 332330
rect 97906 322960 97962 322969
rect 97906 322895 97962 322904
rect 97920 314566 97948 322895
rect 97908 314560 97960 314566
rect 97908 314502 97960 314508
rect 99484 311846 99512 332302
rect 119448 313698 119476 335378
rect 120724 335368 120776 335374
rect 120724 335310 120776 335316
rect 119370 313670 119476 313698
rect 99472 311840 99524 311846
rect 99472 311782 99524 311788
rect 100036 311778 100064 313140
rect 100024 311772 100076 311778
rect 100024 311714 100076 311720
rect 109696 311710 109724 313140
rect 120736 311710 120764 335310
rect 137664 332860 137692 335378
rect 147312 335368 147364 335374
rect 147312 335310 147364 335316
rect 147324 332860 147352 335310
rect 127084 332302 128018 332330
rect 126886 322960 126942 322969
rect 126886 322895 126942 322904
rect 121458 322008 121514 322017
rect 121458 321943 121514 321952
rect 121472 314634 121500 321943
rect 126900 314634 126928 322895
rect 121460 314628 121512 314634
rect 121460 314570 121512 314576
rect 126888 314628 126940 314634
rect 126888 314570 126940 314576
rect 127084 311846 127112 332302
rect 148336 316034 148364 335446
rect 156328 335436 156380 335442
rect 156328 335378 156380 335384
rect 148416 335368 148468 335374
rect 148416 335310 148468 335316
rect 147784 316006 148364 316034
rect 147784 313698 147812 316006
rect 147338 313670 147812 313698
rect 127072 311840 127124 311846
rect 127072 311782 127124 311788
rect 128004 311778 128032 313140
rect 127992 311772 128044 311778
rect 127992 311714 128044 311720
rect 137664 311710 137692 313140
rect 148428 311710 148456 335310
rect 156340 332874 156368 335378
rect 165632 333146 165660 335446
rect 175280 335368 175332 335374
rect 175280 335310 175332 335316
rect 175292 333146 175320 335310
rect 165632 333118 165706 333146
rect 175292 333118 175366 333146
rect 156032 332846 156368 332874
rect 165678 332860 165706 333118
rect 175338 332860 175366 333118
rect 154486 322960 154542 322969
rect 154486 322895 154542 322904
rect 149058 322008 149114 322017
rect 149058 321943 149114 321952
rect 149072 314566 149100 321943
rect 154500 314566 154528 322895
rect 149060 314560 149112 314566
rect 149060 314502 149112 314508
rect 154488 314560 154540 314566
rect 154488 314502 154540 314508
rect 175476 313698 175504 335446
rect 178684 335436 178736 335442
rect 178684 335378 178736 335384
rect 177304 335368 177356 335374
rect 177304 335310 177356 335316
rect 175352 313670 175504 313698
rect 156032 313126 156092 313154
rect 165692 313126 166028 313154
rect 156064 311778 156092 313126
rect 166000 311778 166028 313126
rect 177316 311778 177344 335310
rect 178038 322008 178094 322017
rect 178038 321943 178094 321952
rect 178052 314634 178080 321943
rect 178040 314628 178092 314634
rect 178040 314570 178092 314576
rect 178696 311778 178724 335378
rect 193692 332860 193720 335446
rect 203340 335368 203392 335374
rect 203340 335310 203392 335316
rect 203352 332860 203380 335310
rect 183664 332302 184046 332330
rect 182086 322960 182142 322969
rect 182086 322895 182142 322904
rect 182100 314634 182128 322895
rect 182088 314628 182140 314634
rect 182088 314570 182140 314576
rect 183664 311846 183692 332302
rect 203536 313698 203564 335446
rect 204904 335368 204956 335374
rect 204904 335310 204956 335316
rect 203366 313670 203564 313698
rect 183652 311840 183704 311846
rect 183652 311782 183704 311788
rect 184032 311778 184060 313140
rect 156052 311772 156104 311778
rect 156052 311714 156104 311720
rect 165988 311772 166040 311778
rect 165988 311714 166040 311720
rect 177304 311772 177356 311778
rect 177304 311714 177356 311720
rect 178684 311772 178736 311778
rect 178684 311714 178736 311720
rect 184020 311772 184072 311778
rect 184020 311714 184072 311720
rect 193692 311710 193720 313140
rect 204916 311710 204944 335310
rect 212276 332874 212304 335514
rect 221372 335504 221424 335510
rect 221372 335446 221424 335452
rect 212060 332846 212304 332874
rect 221384 332874 221412 335446
rect 232504 335436 232556 335442
rect 232504 335378 232556 335384
rect 231032 335368 231084 335374
rect 231032 335310 231084 335316
rect 231044 332874 231072 335310
rect 221384 332846 221720 332874
rect 231044 332846 231380 332874
rect 209688 331288 209740 331294
rect 209688 331230 209740 331236
rect 209700 323921 209728 331230
rect 209686 323912 209742 323921
rect 209686 323847 209742 323856
rect 205638 322008 205694 322017
rect 205638 321943 205694 321952
rect 205652 314566 205680 321943
rect 232516 316034 232544 335378
rect 232596 335368 232648 335374
rect 232596 335310 232648 335316
rect 231872 316006 232544 316034
rect 205640 314560 205692 314566
rect 205640 314502 205692 314508
rect 231872 313834 231900 316006
rect 231780 313806 231900 313834
rect 231780 313698 231808 313806
rect 231380 313670 231808 313698
rect 211724 313126 212060 313154
rect 221720 313126 222056 313154
rect 211724 311778 211752 313126
rect 222028 311778 222056 313126
rect 232608 311778 232636 335310
rect 232700 315178 232728 335514
rect 233238 322008 233294 322017
rect 233238 321943 233294 321952
rect 232688 315172 232740 315178
rect 232688 315114 232740 315120
rect 233252 314634 233280 321943
rect 233240 314628 233292 314634
rect 233240 314570 233292 314576
rect 211712 311772 211764 311778
rect 211712 311714 211764 311720
rect 222016 311772 222068 311778
rect 222016 311714 222068 311720
rect 232596 311772 232648 311778
rect 232596 311714 232648 311720
rect 81992 311704 82044 311710
rect 81992 311646 82044 311652
rect 94504 311704 94556 311710
rect 94504 311646 94556 311652
rect 109684 311704 109736 311710
rect 109684 311646 109736 311652
rect 120724 311704 120776 311710
rect 120724 311646 120776 311652
rect 137652 311704 137704 311710
rect 137652 311646 137704 311652
rect 148416 311704 148468 311710
rect 148416 311646 148468 311652
rect 193680 311704 193732 311710
rect 193680 311646 193732 311652
rect 204904 311704 204956 311710
rect 204904 311646 204956 311652
rect 148324 308032 148376 308038
rect 148324 307974 148376 307980
rect 165620 308032 165672 308038
rect 165620 307974 165672 307980
rect 175464 308032 175516 308038
rect 175464 307974 175516 307980
rect 193680 308032 193732 308038
rect 193680 307974 193732 307980
rect 203524 308032 203576 308038
rect 203524 307974 203576 307980
rect 221372 308032 221424 308038
rect 221372 307974 221424 307980
rect 81440 307964 81492 307970
rect 81440 307906 81492 307912
rect 91468 307964 91520 307970
rect 91468 307906 91520 307912
rect 109684 307964 109736 307970
rect 109684 307906 109736 307912
rect 119436 307964 119488 307970
rect 119436 307906 119488 307912
rect 137652 307964 137704 307970
rect 137652 307906 137704 307912
rect 81452 305946 81480 307906
rect 91100 307896 91152 307902
rect 91100 307838 91152 307844
rect 91112 305946 91140 307838
rect 81452 305918 81696 305946
rect 91112 305918 91356 305946
rect 71884 305238 72036 305266
rect 71044 284232 71096 284238
rect 71044 284174 71096 284180
rect 71884 284170 71912 305238
rect 91480 286770 91508 307906
rect 94504 307896 94556 307902
rect 94504 307838 94556 307844
rect 93858 295624 93914 295633
rect 93858 295559 93914 295568
rect 93872 286958 93900 295559
rect 93860 286952 93912 286958
rect 93860 286894 93912 286900
rect 91356 286742 91508 286770
rect 72036 286062 72096 286090
rect 81696 286062 82032 286090
rect 71872 284164 71924 284170
rect 71872 284106 71924 284112
rect 72068 284102 72096 286062
rect 82004 284102 82032 286062
rect 94516 284102 94544 307838
rect 109696 305932 109724 307906
rect 119344 307896 119396 307902
rect 119344 307838 119396 307844
rect 119356 305932 119384 307838
rect 99484 305238 100050 305266
rect 97906 296304 97962 296313
rect 97906 296239 97962 296248
rect 97920 286958 97948 296239
rect 97908 286952 97960 286958
rect 97908 286894 97960 286900
rect 99484 284102 99512 305238
rect 119448 286770 119476 307906
rect 120724 307896 120776 307902
rect 120724 307838 120776 307844
rect 119370 286742 119476 286770
rect 100036 284170 100064 286076
rect 100024 284164 100076 284170
rect 100024 284106 100076 284112
rect 109696 284102 109724 286076
rect 120736 284102 120764 307838
rect 137664 305932 137692 307906
rect 147312 307896 147364 307902
rect 147312 307838 147364 307844
rect 147324 305932 147352 307838
rect 127084 305238 128018 305266
rect 126886 296304 126942 296313
rect 126886 296239 126942 296248
rect 121458 295624 121514 295633
rect 121458 295559 121514 295568
rect 121472 287026 121500 295559
rect 126900 287026 126928 296239
rect 121460 287020 121512 287026
rect 121460 286962 121512 286968
rect 126888 287020 126940 287026
rect 126888 286962 126940 286968
rect 127084 284102 127112 305238
rect 148336 287054 148364 307974
rect 156328 307964 156380 307970
rect 156328 307906 156380 307912
rect 148416 307896 148468 307902
rect 148416 307838 148468 307844
rect 147784 287026 148364 287054
rect 147784 286770 147812 287026
rect 147338 286742 147812 286770
rect 128004 284170 128032 286076
rect 127992 284164 128044 284170
rect 127992 284106 128044 284112
rect 137664 284102 137692 286076
rect 148428 284102 148456 307838
rect 156340 305946 156368 307906
rect 165632 306082 165660 307974
rect 175280 307896 175332 307902
rect 175280 307838 175332 307844
rect 175292 306082 175320 307838
rect 165632 306054 165706 306082
rect 175292 306054 175366 306082
rect 156032 305918 156368 305946
rect 165678 305932 165706 306054
rect 175338 305932 175366 306054
rect 154486 296304 154542 296313
rect 154486 296239 154542 296248
rect 149058 295624 149114 295633
rect 149058 295559 149114 295568
rect 149072 286958 149100 295559
rect 154500 286958 154528 296239
rect 149060 286952 149112 286958
rect 149060 286894 149112 286900
rect 154488 286952 154540 286958
rect 154488 286894 154540 286900
rect 175476 286770 175504 307974
rect 178684 307964 178736 307970
rect 178684 307906 178736 307912
rect 177304 307896 177356 307902
rect 177304 307838 177356 307844
rect 175352 286742 175504 286770
rect 156032 286062 156092 286090
rect 165692 286062 166028 286090
rect 156064 284170 156092 286062
rect 166000 284170 166028 286062
rect 177316 284170 177344 307838
rect 178038 295624 178094 295633
rect 178038 295559 178094 295568
rect 178052 287026 178080 295559
rect 178040 287020 178092 287026
rect 178040 286962 178092 286968
rect 178696 284306 178724 307906
rect 193692 305932 193720 307974
rect 203340 307896 203392 307902
rect 203340 307838 203392 307844
rect 203352 305932 203380 307838
rect 183664 305238 184046 305266
rect 182086 296304 182142 296313
rect 182086 296239 182142 296248
rect 182100 286890 182128 296239
rect 182088 286884 182140 286890
rect 182088 286826 182140 286832
rect 178684 284300 178736 284306
rect 178684 284242 178736 284248
rect 183664 284170 183692 305238
rect 203536 286770 203564 307974
rect 204904 307896 204956 307902
rect 204904 307838 204956 307844
rect 203366 286742 203564 286770
rect 184032 284306 184060 286076
rect 184020 284300 184072 284306
rect 184020 284242 184072 284248
rect 156052 284164 156104 284170
rect 156052 284106 156104 284112
rect 165988 284164 166040 284170
rect 165988 284106 166040 284112
rect 177304 284164 177356 284170
rect 177304 284106 177356 284112
rect 183652 284164 183704 284170
rect 183652 284106 183704 284112
rect 193692 284102 193720 286076
rect 204916 284102 204944 307838
rect 212264 307828 212316 307834
rect 212264 307770 212316 307776
rect 212276 305946 212304 307770
rect 212060 305918 212304 305946
rect 221384 305946 221412 307974
rect 232596 307964 232648 307970
rect 232596 307906 232648 307912
rect 231032 307896 231084 307902
rect 231032 307838 231084 307844
rect 232504 307896 232556 307902
rect 232504 307838 232556 307844
rect 231044 305946 231072 307838
rect 221384 305918 221720 305946
rect 231044 305918 231380 305946
rect 209686 296304 209742 296313
rect 209686 296239 209742 296248
rect 205638 295624 205694 295633
rect 205638 295559 205694 295568
rect 205652 286958 205680 295559
rect 209700 287026 209728 296239
rect 209688 287020 209740 287026
rect 209688 286962 209740 286968
rect 205640 286952 205692 286958
rect 205640 286894 205692 286900
rect 231676 286816 231728 286822
rect 231380 286764 231676 286770
rect 231380 286758 231728 286764
rect 231380 286742 231716 286758
rect 211724 286062 212060 286090
rect 221720 286062 222056 286090
rect 211724 284170 211752 286062
rect 222028 284170 222056 286062
rect 232516 284170 232544 307838
rect 232608 286822 232636 307906
rect 232688 307828 232740 307834
rect 232688 307770 232740 307776
rect 232700 287978 232728 307770
rect 233238 295624 233294 295633
rect 233238 295559 233294 295568
rect 232688 287972 232740 287978
rect 232688 287914 232740 287920
rect 233252 286890 233280 295559
rect 233240 286884 233292 286890
rect 233240 286826 233292 286832
rect 232596 286816 232648 286822
rect 232596 286758 232648 286764
rect 211712 284164 211764 284170
rect 211712 284106 211764 284112
rect 222016 284164 222068 284170
rect 222016 284106 222068 284112
rect 232504 284164 232556 284170
rect 232504 284106 232556 284112
rect 72056 284096 72108 284102
rect 72056 284038 72108 284044
rect 81992 284096 82044 284102
rect 81992 284038 82044 284044
rect 94504 284096 94556 284102
rect 94504 284038 94556 284044
rect 99472 284096 99524 284102
rect 99472 284038 99524 284044
rect 109684 284096 109736 284102
rect 109684 284038 109736 284044
rect 120724 284096 120776 284102
rect 120724 284038 120776 284044
rect 127072 284096 127124 284102
rect 127072 284038 127124 284044
rect 137652 284096 137704 284102
rect 137652 284038 137704 284044
rect 148416 284096 148468 284102
rect 148416 284038 148468 284044
rect 193680 284096 193732 284102
rect 193680 284038 193732 284044
rect 204904 284096 204956 284102
rect 204904 284038 204956 284044
rect 71044 280424 71096 280430
rect 71044 280366 71096 280372
rect 212356 280424 212408 280430
rect 212356 280366 212408 280372
rect 232688 280424 232740 280430
rect 232688 280366 232740 280372
rect 69664 280220 69716 280226
rect 69664 280162 69716 280168
rect 69676 256562 69704 280162
rect 70308 277432 70360 277438
rect 70308 277374 70360 277380
rect 70320 269793 70348 277374
rect 70306 269784 70362 269793
rect 70306 269719 70362 269728
rect 69664 256556 69716 256562
rect 69664 256498 69716 256504
rect 69664 254176 69716 254182
rect 69664 254118 69716 254124
rect 69676 202774 69704 254118
rect 70306 242312 70362 242321
rect 70306 242247 70362 242256
rect 70320 233238 70348 242247
rect 70308 233232 70360 233238
rect 70308 233174 70360 233180
rect 71056 230382 71084 280366
rect 148416 280356 148468 280362
rect 148416 280298 148468 280304
rect 165712 280356 165764 280362
rect 165712 280298 165764 280304
rect 175464 280356 175516 280362
rect 175464 280298 175516 280304
rect 193680 280356 193732 280362
rect 193680 280298 193732 280304
rect 203524 280356 203576 280362
rect 203524 280298 203576 280304
rect 81440 280288 81492 280294
rect 81440 280230 81492 280236
rect 91468 280288 91520 280294
rect 91468 280230 91520 280236
rect 109684 280288 109736 280294
rect 109684 280230 109736 280236
rect 119436 280288 119488 280294
rect 119436 280230 119488 280236
rect 137652 280288 137704 280294
rect 137652 280230 137704 280236
rect 81452 278882 81480 280230
rect 91100 280220 91152 280226
rect 91100 280162 91152 280168
rect 91112 278882 91140 280162
rect 81452 278854 81696 278882
rect 91112 278854 91356 278882
rect 71884 278310 72036 278338
rect 71884 256630 71912 278310
rect 91480 259706 91508 280230
rect 94504 280220 94556 280226
rect 94504 280162 94556 280168
rect 93860 277500 93912 277506
rect 93860 277442 93912 277448
rect 93872 268569 93900 277442
rect 93858 268560 93914 268569
rect 93858 268495 93914 268504
rect 91356 259678 91508 259706
rect 72022 258890 72050 259148
rect 81696 259134 82032 259162
rect 71976 258862 72050 258890
rect 71976 256698 72004 258862
rect 71964 256692 72016 256698
rect 71964 256634 72016 256640
rect 71872 256624 71924 256630
rect 71872 256566 71924 256572
rect 82004 256562 82032 259134
rect 94516 256562 94544 280162
rect 109696 278868 109724 280230
rect 119344 280220 119396 280226
rect 119344 280162 119396 280168
rect 119356 278868 119384 280162
rect 99484 278310 100050 278338
rect 97908 277500 97960 277506
rect 97908 277442 97960 277448
rect 97920 269249 97948 277442
rect 97906 269240 97962 269249
rect 97906 269175 97962 269184
rect 99484 256698 99512 278310
rect 119448 259706 119476 280230
rect 120724 280220 120776 280226
rect 120724 280162 120776 280168
rect 119370 259678 119476 259706
rect 99472 256692 99524 256698
rect 99472 256634 99524 256640
rect 100036 256630 100064 259148
rect 100024 256624 100076 256630
rect 100024 256566 100076 256572
rect 109696 256562 109724 259148
rect 120736 256562 120764 280162
rect 137664 278868 137692 280230
rect 147312 280220 147364 280226
rect 147312 280162 147364 280168
rect 148324 280220 148376 280226
rect 148324 280162 148376 280168
rect 147324 278868 147352 280162
rect 127084 278310 128018 278338
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 126888 277432 126940 277438
rect 126888 277374 126940 277380
rect 121472 268569 121500 277374
rect 126900 269249 126928 277374
rect 126886 269240 126942 269249
rect 126886 269175 126942 269184
rect 121458 268560 121514 268569
rect 121458 268495 121514 268504
rect 127084 256698 127112 278310
rect 147680 259480 147732 259486
rect 147338 259428 147680 259434
rect 147338 259422 147732 259428
rect 147338 259406 147720 259422
rect 127072 256692 127124 256698
rect 127072 256634 127124 256640
rect 128004 256630 128032 259148
rect 127992 256624 128044 256630
rect 127992 256566 128044 256572
rect 137664 256562 137692 259148
rect 148336 256562 148364 280162
rect 148428 259486 148456 280298
rect 156328 280288 156380 280294
rect 156328 280230 156380 280236
rect 156340 278882 156368 280230
rect 156032 278854 156368 278882
rect 165724 278746 165752 280298
rect 175372 280220 175424 280226
rect 175372 280162 175424 280168
rect 175384 278746 175412 280162
rect 165692 278718 165752 278746
rect 175352 278718 175412 278746
rect 149060 277500 149112 277506
rect 149060 277442 149112 277448
rect 154488 277500 154540 277506
rect 154488 277442 154540 277448
rect 149072 268569 149100 277442
rect 154500 269249 154528 277442
rect 154486 269240 154542 269249
rect 154486 269175 154542 269184
rect 149058 268560 149114 268569
rect 149058 268495 149114 268504
rect 175476 259706 175504 280298
rect 178684 280288 178736 280294
rect 178684 280230 178736 280236
rect 177304 280220 177356 280226
rect 177304 280162 177356 280168
rect 175352 259678 175504 259706
rect 148416 259480 148468 259486
rect 148416 259422 148468 259428
rect 156018 258890 156046 259148
rect 165692 259134 166028 259162
rect 155972 258862 156046 258890
rect 155972 256630 156000 258862
rect 166000 256630 166028 259134
rect 177316 256630 177344 280162
rect 178040 277432 178092 277438
rect 178040 277374 178092 277380
rect 178052 268569 178080 277374
rect 178038 268560 178094 268569
rect 178038 268495 178094 268504
rect 178696 256630 178724 280230
rect 193692 278868 193720 280298
rect 203340 280220 203392 280226
rect 203340 280162 203392 280168
rect 203352 278868 203380 280162
rect 183664 278310 184046 278338
rect 182088 277568 182140 277574
rect 182088 277510 182140 277516
rect 182100 269249 182128 277510
rect 182086 269240 182142 269249
rect 182086 269175 182142 269184
rect 183664 256698 183692 278310
rect 203536 259706 203564 280298
rect 204904 280220 204956 280226
rect 204904 280162 204956 280168
rect 203366 259678 203564 259706
rect 183652 256692 183704 256698
rect 183652 256634 183704 256640
rect 184032 256630 184060 259148
rect 155960 256624 156012 256630
rect 155960 256566 156012 256572
rect 165988 256624 166040 256630
rect 165988 256566 166040 256572
rect 177304 256624 177356 256630
rect 177304 256566 177356 256572
rect 178684 256624 178736 256630
rect 178684 256566 178736 256572
rect 184020 256624 184072 256630
rect 184020 256566 184072 256572
rect 193692 256562 193720 259148
rect 204916 256562 204944 280162
rect 212368 278882 212396 280366
rect 221372 280356 221424 280362
rect 221372 280298 221424 280304
rect 212060 278854 212396 278882
rect 221384 278882 221412 280298
rect 232504 280288 232556 280294
rect 232504 280230 232556 280236
rect 231032 280220 231084 280226
rect 231032 280162 231084 280168
rect 231044 278882 231072 280162
rect 221384 278854 221720 278882
rect 231044 278854 231380 278882
rect 205640 277500 205692 277506
rect 205640 277442 205692 277448
rect 205652 269113 205680 277442
rect 209688 277432 209740 277438
rect 209688 277374 209740 277380
rect 209700 269249 209728 277374
rect 209686 269240 209742 269249
rect 209686 269175 209742 269184
rect 205638 269104 205694 269113
rect 205638 269039 205694 269048
rect 232516 267734 232544 280230
rect 232596 280220 232648 280226
rect 232596 280162 232648 280168
rect 231872 267706 232544 267734
rect 231872 259434 231900 267706
rect 231380 259406 231900 259434
rect 211724 259134 212060 259162
rect 221720 259134 221964 259162
rect 211724 256630 211752 259134
rect 221936 256630 221964 259134
rect 232608 256630 232636 280162
rect 232700 262206 232728 280366
rect 233240 277568 233292 277574
rect 233240 277510 233292 277516
rect 233252 268569 233280 277510
rect 233238 268560 233294 268569
rect 233238 268495 233294 268504
rect 232688 262200 232740 262206
rect 232688 262142 232740 262148
rect 211712 256624 211764 256630
rect 211712 256566 211764 256572
rect 221924 256624 221976 256630
rect 221924 256566 221976 256572
rect 232596 256624 232648 256630
rect 232596 256566 232648 256572
rect 81992 256556 82044 256562
rect 81992 256498 82044 256504
rect 94504 256556 94556 256562
rect 94504 256498 94556 256504
rect 109684 256556 109736 256562
rect 109684 256498 109736 256504
rect 120724 256556 120776 256562
rect 120724 256498 120776 256504
rect 137652 256556 137704 256562
rect 137652 256498 137704 256504
rect 148324 256556 148376 256562
rect 148324 256498 148376 256504
rect 193680 256556 193732 256562
rect 193680 256498 193732 256504
rect 204904 256556 204956 256562
rect 204904 256498 204956 256504
rect 212356 254176 212408 254182
rect 212356 254118 212408 254124
rect 232688 254176 232740 254182
rect 232688 254118 232740 254124
rect 81440 254108 81492 254114
rect 81440 254050 81492 254056
rect 148416 254108 148468 254114
rect 148416 254050 148468 254056
rect 165712 254108 165764 254114
rect 165712 254050 165764 254056
rect 175464 254108 175516 254114
rect 175464 254050 175516 254056
rect 193680 254108 193732 254114
rect 193680 254050 193732 254056
rect 203524 254108 203576 254114
rect 203524 254050 203576 254056
rect 81452 251954 81480 254050
rect 91100 254040 91152 254046
rect 91100 253982 91152 253988
rect 91468 254040 91520 254046
rect 91468 253982 91520 253988
rect 109684 254040 109736 254046
rect 109684 253982 109736 253988
rect 119436 254040 119488 254046
rect 119436 253982 119488 253988
rect 137652 254040 137704 254046
rect 137652 253982 137704 253988
rect 91112 251954 91140 253982
rect 81452 251926 81696 251954
rect 91112 251926 91356 251954
rect 71884 251246 72036 251274
rect 71044 230376 71096 230382
rect 71044 230318 71096 230324
rect 71884 230314 71912 251246
rect 91480 232778 91508 253982
rect 94504 253972 94556 253978
rect 94504 253914 94556 253920
rect 93860 251252 93912 251258
rect 93860 251194 93912 251200
rect 93872 241641 93900 251194
rect 93858 241632 93914 241641
rect 93858 241567 93914 241576
rect 91356 232750 91508 232778
rect 72036 232070 72096 232098
rect 81696 232070 82032 232098
rect 71872 230308 71924 230314
rect 71872 230250 71924 230256
rect 72068 230246 72096 232070
rect 82004 230246 82032 232070
rect 94516 230246 94544 253914
rect 109696 251940 109724 253982
rect 119344 253972 119396 253978
rect 119344 253914 119396 253920
rect 119356 251940 119384 253914
rect 97908 251252 97960 251258
rect 97908 251194 97960 251200
rect 99484 251246 100050 251274
rect 97920 242321 97948 251194
rect 97906 242312 97962 242321
rect 97906 242247 97962 242256
rect 99484 230246 99512 251246
rect 119448 232778 119476 253982
rect 120724 253972 120776 253978
rect 120724 253914 120776 253920
rect 119370 232750 119476 232778
rect 100036 230314 100064 232084
rect 100024 230308 100076 230314
rect 100024 230250 100076 230256
rect 109696 230246 109724 232084
rect 120736 230246 120764 253914
rect 137664 251940 137692 253982
rect 147312 253972 147364 253978
rect 147312 253914 147364 253920
rect 148324 253972 148376 253978
rect 148324 253914 148376 253920
rect 147324 251940 147352 253914
rect 127084 251246 128018 251274
rect 126886 242312 126942 242321
rect 126886 242247 126942 242256
rect 121458 241632 121514 241641
rect 121458 241567 121514 241576
rect 121472 233238 121500 241567
rect 126900 233238 126928 242247
rect 121460 233232 121512 233238
rect 121460 233174 121512 233180
rect 126888 233232 126940 233238
rect 126888 233174 126940 233180
rect 127084 230246 127112 251246
rect 147680 235408 147732 235414
rect 147680 235350 147732 235356
rect 147692 232778 147720 235350
rect 147338 232750 147720 232778
rect 128004 230314 128032 232084
rect 127992 230308 128044 230314
rect 127992 230250 128044 230256
rect 137664 230246 137692 232084
rect 148336 230246 148364 253914
rect 148428 235414 148456 254050
rect 156328 254040 156380 254046
rect 156328 253982 156380 253988
rect 156340 251954 156368 253982
rect 156032 251926 156368 251954
rect 165724 251818 165752 254050
rect 175372 253972 175424 253978
rect 175372 253914 175424 253920
rect 175384 251818 175412 253914
rect 165692 251790 165752 251818
rect 175352 251790 175412 251818
rect 149060 251252 149112 251258
rect 149060 251194 149112 251200
rect 154488 251252 154540 251258
rect 154488 251194 154540 251200
rect 149072 241641 149100 251194
rect 154500 242321 154528 251194
rect 154486 242312 154542 242321
rect 154486 242247 154542 242256
rect 149058 241632 149114 241641
rect 149058 241567 149114 241576
rect 148416 235408 148468 235414
rect 148416 235350 148468 235356
rect 175476 232778 175504 254050
rect 178684 254040 178736 254046
rect 178684 253982 178736 253988
rect 177304 253972 177356 253978
rect 177304 253914 177356 253920
rect 175352 232750 175504 232778
rect 156032 232070 156092 232098
rect 165692 232070 166028 232098
rect 156064 230314 156092 232070
rect 166000 230314 166028 232070
rect 177316 230314 177344 253914
rect 178038 241632 178094 241641
rect 178038 241567 178094 241576
rect 178052 233238 178080 241567
rect 178040 233232 178092 233238
rect 178040 233174 178092 233180
rect 178696 230450 178724 253982
rect 193692 251940 193720 254050
rect 203340 253972 203392 253978
rect 203340 253914 203392 253920
rect 203352 251940 203380 253914
rect 182088 251320 182140 251326
rect 182088 251262 182140 251268
rect 182100 242321 182128 251262
rect 183664 251246 184046 251274
rect 182086 242312 182142 242321
rect 182086 242247 182142 242256
rect 178684 230444 178736 230450
rect 178684 230386 178736 230392
rect 183664 230314 183692 251246
rect 203536 232778 203564 254050
rect 204904 253972 204956 253978
rect 204904 253914 204956 253920
rect 203366 232750 203564 232778
rect 184032 230450 184060 232084
rect 184020 230444 184072 230450
rect 184020 230386 184072 230392
rect 156052 230308 156104 230314
rect 156052 230250 156104 230256
rect 165988 230308 166040 230314
rect 165988 230250 166040 230256
rect 177304 230308 177356 230314
rect 177304 230250 177356 230256
rect 183652 230308 183704 230314
rect 183652 230250 183704 230256
rect 193692 230246 193720 232084
rect 204916 230246 204944 253914
rect 212368 251954 212396 254118
rect 221372 254108 221424 254114
rect 221372 254050 221424 254056
rect 212060 251926 212396 251954
rect 221384 251954 221412 254050
rect 232596 254040 232648 254046
rect 232596 253982 232648 253988
rect 231032 253972 231084 253978
rect 231032 253914 231084 253920
rect 232504 253972 232556 253978
rect 232504 253914 232556 253920
rect 231044 251954 231072 253914
rect 221384 251926 221720 251954
rect 231044 251926 231380 251954
rect 205640 251252 205692 251258
rect 205640 251194 205692 251200
rect 205652 241641 205680 251194
rect 209686 242312 209742 242321
rect 209686 242247 209742 242256
rect 205638 241632 205694 241641
rect 205638 241567 205694 241576
rect 209700 233238 209728 242247
rect 209688 233232 209740 233238
rect 209688 233174 209740 233180
rect 231676 233164 231728 233170
rect 231676 233106 231728 233112
rect 231688 232778 231716 233106
rect 231380 232750 231716 232778
rect 211724 232070 212060 232098
rect 221720 232070 222056 232098
rect 211724 230314 211752 232070
rect 222028 230314 222056 232070
rect 232516 230314 232544 253914
rect 232608 233170 232636 253982
rect 232700 233578 232728 254118
rect 233240 251320 233292 251326
rect 233240 251262 233292 251268
rect 233252 241641 233280 251262
rect 233238 241632 233294 241641
rect 233238 241567 233294 241576
rect 232688 233572 232740 233578
rect 232688 233514 232740 233520
rect 232596 233164 232648 233170
rect 232596 233106 232648 233112
rect 211712 230308 211764 230314
rect 211712 230250 211764 230256
rect 222016 230308 222068 230314
rect 222016 230250 222068 230256
rect 232504 230308 232556 230314
rect 232504 230250 232556 230256
rect 72056 230240 72108 230246
rect 72056 230182 72108 230188
rect 81992 230240 82044 230246
rect 81992 230182 82044 230188
rect 94504 230240 94556 230246
rect 94504 230182 94556 230188
rect 99472 230240 99524 230246
rect 99472 230182 99524 230188
rect 109684 230240 109736 230246
rect 109684 230182 109736 230188
rect 120724 230240 120776 230246
rect 120724 230182 120776 230188
rect 127072 230240 127124 230246
rect 127072 230182 127124 230188
rect 137652 230240 137704 230246
rect 137652 230182 137704 230188
rect 148324 230240 148376 230246
rect 148324 230182 148376 230188
rect 193680 230240 193732 230246
rect 193680 230182 193732 230188
rect 204904 230240 204956 230246
rect 204904 230182 204956 230188
rect 148324 226568 148376 226574
rect 148324 226510 148376 226516
rect 165712 226568 165764 226574
rect 165712 226510 165764 226516
rect 175464 226568 175516 226574
rect 175464 226510 175516 226516
rect 193680 226568 193732 226574
rect 193680 226510 193732 226516
rect 203524 226568 203576 226574
rect 203524 226510 203576 226516
rect 221372 226568 221424 226574
rect 221372 226510 221424 226516
rect 81440 226500 81492 226506
rect 81440 226442 81492 226448
rect 91468 226500 91520 226506
rect 91468 226442 91520 226448
rect 109684 226500 109736 226506
rect 109684 226442 109736 226448
rect 119436 226500 119488 226506
rect 119436 226442 119488 226448
rect 137652 226500 137704 226506
rect 137652 226442 137704 226448
rect 81452 224890 81480 226442
rect 91100 226432 91152 226438
rect 91100 226374 91152 226380
rect 91112 224890 91140 226374
rect 81452 224862 81696 224890
rect 91112 224862 91356 224890
rect 71884 224318 72036 224346
rect 70306 214704 70362 214713
rect 70306 214639 70362 214648
rect 70320 205630 70348 214639
rect 70308 205624 70360 205630
rect 70308 205566 70360 205572
rect 69664 202768 69716 202774
rect 69664 202710 69716 202716
rect 71884 202706 71912 224318
rect 91480 205714 91508 226442
rect 94504 226432 94556 226438
rect 94504 226374 94556 226380
rect 93858 214568 93914 214577
rect 93858 214503 93914 214512
rect 91356 205686 91508 205714
rect 93872 205562 93900 214503
rect 93860 205556 93912 205562
rect 93860 205498 93912 205504
rect 72036 205006 72096 205034
rect 81696 205006 82032 205034
rect 71872 202700 71924 202706
rect 71872 202642 71924 202648
rect 72068 202638 72096 205006
rect 82004 202638 82032 205006
rect 94516 202638 94544 226374
rect 109696 224876 109724 226442
rect 119344 226432 119396 226438
rect 119344 226374 119396 226380
rect 119356 224876 119384 226374
rect 99484 224318 100050 224346
rect 97906 215248 97962 215257
rect 97906 215183 97962 215192
rect 97920 205562 97948 215183
rect 97908 205556 97960 205562
rect 97908 205498 97960 205504
rect 99484 202638 99512 224318
rect 119448 205714 119476 226442
rect 120724 226432 120776 226438
rect 120724 226374 120776 226380
rect 119370 205686 119476 205714
rect 100036 202706 100064 205020
rect 100024 202700 100076 202706
rect 100024 202642 100076 202648
rect 109696 202638 109724 205020
rect 120736 202638 120764 226374
rect 137664 224876 137692 226442
rect 147312 226432 147364 226438
rect 147312 226374 147364 226380
rect 147324 224876 147352 226374
rect 127084 224318 128018 224346
rect 126886 215248 126942 215257
rect 126886 215183 126942 215192
rect 121458 214568 121514 214577
rect 121458 214503 121514 214512
rect 121472 205630 121500 214503
rect 126900 205630 126928 215183
rect 121460 205624 121512 205630
rect 121460 205566 121512 205572
rect 126888 205624 126940 205630
rect 126888 205566 126940 205572
rect 127084 202638 127112 224318
rect 148336 209774 148364 226510
rect 156328 226500 156380 226506
rect 156328 226442 156380 226448
rect 148416 226432 148468 226438
rect 148416 226374 148468 226380
rect 147784 209746 148364 209774
rect 147784 205578 147812 209746
rect 147338 205550 147812 205578
rect 127728 205006 128018 205034
rect 137678 205006 137968 205034
rect 127728 202706 127756 205006
rect 127716 202700 127768 202706
rect 127716 202642 127768 202648
rect 137940 202638 137968 205006
rect 148428 202638 148456 226374
rect 156340 224890 156368 226442
rect 156032 224862 156368 224890
rect 165724 224754 165752 226510
rect 175372 226432 175424 226438
rect 175372 226374 175424 226380
rect 175384 224754 175412 226374
rect 165692 224726 165752 224754
rect 175352 224726 175412 224754
rect 154486 215248 154542 215257
rect 154486 215183 154542 215192
rect 149058 214568 149114 214577
rect 149058 214503 149114 214512
rect 149072 205562 149100 214503
rect 154500 205562 154528 215183
rect 175476 205714 175504 226510
rect 178684 226500 178736 226506
rect 178684 226442 178736 226448
rect 177304 226432 177356 226438
rect 177304 226374 177356 226380
rect 175352 205686 175504 205714
rect 149060 205556 149112 205562
rect 149060 205498 149112 205504
rect 154488 205556 154540 205562
rect 154488 205498 154540 205504
rect 156032 205006 156092 205034
rect 165692 205006 166028 205034
rect 156064 202706 156092 205006
rect 166000 202706 166028 205006
rect 177316 202706 177344 226374
rect 178038 214568 178094 214577
rect 178038 214503 178094 214512
rect 178052 205630 178080 214503
rect 178040 205624 178092 205630
rect 178040 205566 178092 205572
rect 178696 202842 178724 226442
rect 193692 224876 193720 226510
rect 203340 226432 203392 226438
rect 203340 226374 203392 226380
rect 203352 224876 203380 226374
rect 183664 224318 184046 224346
rect 182086 215248 182142 215257
rect 182086 215183 182142 215192
rect 182100 205494 182128 215183
rect 182088 205488 182140 205494
rect 182088 205430 182140 205436
rect 178684 202836 178736 202842
rect 178684 202778 178736 202784
rect 183664 202706 183692 224318
rect 203536 205714 203564 226510
rect 204904 226432 204956 226438
rect 204904 226374 204956 226380
rect 203366 205686 203564 205714
rect 184032 202842 184060 205020
rect 184020 202836 184072 202842
rect 184020 202778 184072 202784
rect 156052 202700 156104 202706
rect 156052 202642 156104 202648
rect 165988 202700 166040 202706
rect 165988 202642 166040 202648
rect 177304 202700 177356 202706
rect 177304 202642 177356 202648
rect 183652 202700 183704 202706
rect 183652 202642 183704 202648
rect 193692 202638 193720 205020
rect 204916 202638 204944 226374
rect 212356 226364 212408 226370
rect 212356 226306 212408 226312
rect 212368 224890 212396 226306
rect 212060 224862 212396 224890
rect 221384 224890 221412 226510
rect 232504 226500 232556 226506
rect 232504 226442 232556 226448
rect 231032 226432 231084 226438
rect 231032 226374 231084 226380
rect 231044 224890 231072 226374
rect 221384 224862 221720 224890
rect 231044 224862 231380 224890
rect 209686 215248 209742 215257
rect 209686 215183 209742 215192
rect 205638 214024 205694 214033
rect 205638 213959 205694 213968
rect 205652 205562 205680 213959
rect 209700 205630 209728 215183
rect 232516 209774 232544 226442
rect 232596 226432 232648 226438
rect 232596 226374 232648 226380
rect 231872 209746 232544 209774
rect 209688 205624 209740 205630
rect 231872 205578 231900 209746
rect 209688 205566 209740 205572
rect 205640 205556 205692 205562
rect 231380 205550 231900 205578
rect 205640 205498 205692 205504
rect 211724 205006 212060 205034
rect 221720 205006 222056 205034
rect 211724 202706 211752 205006
rect 222028 202706 222056 205006
rect 232608 202706 232636 226374
rect 232688 226364 232740 226370
rect 232688 226306 232740 226312
rect 232700 207806 232728 226306
rect 233238 214568 233294 214577
rect 233238 214503 233294 214512
rect 232688 207800 232740 207806
rect 232688 207742 232740 207748
rect 233252 205494 233280 214503
rect 233240 205488 233292 205494
rect 233240 205430 233292 205436
rect 211712 202700 211764 202706
rect 211712 202642 211764 202648
rect 222016 202700 222068 202706
rect 222016 202642 222068 202648
rect 232596 202700 232648 202706
rect 232596 202642 232648 202648
rect 72056 202632 72108 202638
rect 72056 202574 72108 202580
rect 81992 202632 82044 202638
rect 81992 202574 82044 202580
rect 94504 202632 94556 202638
rect 94504 202574 94556 202580
rect 99472 202632 99524 202638
rect 99472 202574 99524 202580
rect 109684 202632 109736 202638
rect 109684 202574 109736 202580
rect 120724 202632 120776 202638
rect 120724 202574 120776 202580
rect 127072 202632 127124 202638
rect 127072 202574 127124 202580
rect 137928 202632 137980 202638
rect 137928 202574 137980 202580
rect 148416 202632 148468 202638
rect 148416 202574 148468 202580
rect 193680 202632 193732 202638
rect 193680 202574 193732 202580
rect 204904 202632 204956 202638
rect 204904 202574 204956 202580
rect 71044 200388 71096 200394
rect 71044 200330 71096 200336
rect 212264 200388 212316 200394
rect 212264 200330 212316 200336
rect 232688 200388 232740 200394
rect 232688 200330 232740 200336
rect 69664 200184 69716 200190
rect 69664 200126 69716 200132
rect 69676 176526 69704 200126
rect 70306 188320 70362 188329
rect 70306 188255 70362 188264
rect 70320 179382 70348 188255
rect 70308 179376 70360 179382
rect 70308 179318 70360 179324
rect 69664 176520 69716 176526
rect 69664 176462 69716 176468
rect 70306 161256 70362 161265
rect 70306 161191 70362 161200
rect 70320 151774 70348 161191
rect 70308 151768 70360 151774
rect 70308 151710 70360 151716
rect 71056 148986 71084 200330
rect 148416 200320 148468 200326
rect 148416 200262 148468 200268
rect 165620 200320 165672 200326
rect 165620 200262 165672 200268
rect 175464 200320 175516 200326
rect 175464 200262 175516 200268
rect 193680 200320 193732 200326
rect 193680 200262 193732 200268
rect 203524 200320 203576 200326
rect 203524 200262 203576 200268
rect 81440 200252 81492 200258
rect 81440 200194 81492 200200
rect 91468 200252 91520 200258
rect 91468 200194 91520 200200
rect 109684 200252 109736 200258
rect 109684 200194 109736 200200
rect 119436 200252 119488 200258
rect 119436 200194 119488 200200
rect 137652 200252 137704 200258
rect 137652 200194 137704 200200
rect 81452 197962 81480 200194
rect 91100 200184 91152 200190
rect 91100 200126 91152 200132
rect 91112 197962 91140 200126
rect 81452 197934 81696 197962
rect 91112 197934 91356 197962
rect 71884 197254 72036 197282
rect 71884 176594 71912 197254
rect 91480 178786 91508 200194
rect 94504 200184 94556 200190
rect 94504 200126 94556 200132
rect 93858 187640 93914 187649
rect 93858 187575 93914 187584
rect 93872 179314 93900 187575
rect 93860 179308 93912 179314
rect 93860 179250 93912 179256
rect 91356 178758 91508 178786
rect 72036 178078 72096 178106
rect 81696 178078 82032 178106
rect 72068 176662 72096 178078
rect 72056 176656 72108 176662
rect 72056 176598 72108 176604
rect 71872 176588 71924 176594
rect 71872 176530 71924 176536
rect 82004 176526 82032 178078
rect 94516 176526 94544 200126
rect 109696 197948 109724 200194
rect 119344 200184 119396 200190
rect 119344 200126 119396 200132
rect 119356 197948 119384 200126
rect 99484 197254 100050 197282
rect 97906 188320 97962 188329
rect 97906 188255 97962 188264
rect 97920 179314 97948 188255
rect 97908 179308 97960 179314
rect 97908 179250 97960 179256
rect 99484 176662 99512 197254
rect 119448 178786 119476 200194
rect 120724 200184 120776 200190
rect 120724 200126 120776 200132
rect 119370 178758 119476 178786
rect 99472 176656 99524 176662
rect 99472 176598 99524 176604
rect 100036 176594 100064 178092
rect 100024 176588 100076 176594
rect 100024 176530 100076 176536
rect 109696 176526 109724 178092
rect 120736 176526 120764 200126
rect 137664 197948 137692 200194
rect 147312 200184 147364 200190
rect 147312 200126 147364 200132
rect 148324 200184 148376 200190
rect 148324 200126 148376 200132
rect 147324 197948 147352 200126
rect 127084 197254 128018 197282
rect 126886 188320 126942 188329
rect 126886 188255 126942 188264
rect 121458 187640 121514 187649
rect 121458 187575 121514 187584
rect 121472 179382 121500 187575
rect 126900 179382 126928 188255
rect 121460 179376 121512 179382
rect 121460 179318 121512 179324
rect 126888 179376 126940 179382
rect 126888 179318 126940 179324
rect 127084 176662 127112 197254
rect 147680 185632 147732 185638
rect 147680 185574 147732 185580
rect 147692 178786 147720 185574
rect 147338 178758 147720 178786
rect 127072 176656 127124 176662
rect 127072 176598 127124 176604
rect 128004 176594 128032 178092
rect 127992 176588 128044 176594
rect 127992 176530 128044 176536
rect 137664 176526 137692 178092
rect 148336 176526 148364 200126
rect 148428 185638 148456 200262
rect 156328 200252 156380 200258
rect 156328 200194 156380 200200
rect 156340 197962 156368 200194
rect 165632 198234 165660 200262
rect 175280 200184 175332 200190
rect 175280 200126 175332 200132
rect 175292 198234 175320 200126
rect 165632 198206 165706 198234
rect 175292 198206 175366 198234
rect 156032 197934 156368 197962
rect 165678 197948 165706 198206
rect 175338 197948 175366 198206
rect 154486 188320 154542 188329
rect 154486 188255 154542 188264
rect 149058 187640 149114 187649
rect 149058 187575 149114 187584
rect 148416 185632 148468 185638
rect 148416 185574 148468 185580
rect 149072 179314 149100 187575
rect 154500 179314 154528 188255
rect 149060 179308 149112 179314
rect 149060 179250 149112 179256
rect 154488 179308 154540 179314
rect 154488 179250 154540 179256
rect 175476 178786 175504 200262
rect 178684 200252 178736 200258
rect 178684 200194 178736 200200
rect 177304 200184 177356 200190
rect 177304 200126 177356 200132
rect 175352 178758 175504 178786
rect 156032 178078 156092 178106
rect 165692 178078 166028 178106
rect 156064 176594 156092 178078
rect 166000 176594 166028 178078
rect 177316 176594 177344 200126
rect 178038 187640 178094 187649
rect 178038 187575 178094 187584
rect 178052 179382 178080 187575
rect 178040 179376 178092 179382
rect 178040 179318 178092 179324
rect 178696 176594 178724 200194
rect 193692 197948 193720 200262
rect 203340 200184 203392 200190
rect 203340 200126 203392 200132
rect 203352 197948 203380 200126
rect 183664 197254 184046 197282
rect 182086 188320 182142 188329
rect 182086 188255 182142 188264
rect 182100 179246 182128 188255
rect 182088 179240 182140 179246
rect 182088 179182 182140 179188
rect 183664 176662 183692 197254
rect 203536 178786 203564 200262
rect 204904 200184 204956 200190
rect 204904 200126 204956 200132
rect 203366 178758 203564 178786
rect 183652 176656 183704 176662
rect 183652 176598 183704 176604
rect 184032 176594 184060 178092
rect 156052 176588 156104 176594
rect 156052 176530 156104 176536
rect 165988 176588 166040 176594
rect 165988 176530 166040 176536
rect 177304 176588 177356 176594
rect 177304 176530 177356 176536
rect 178684 176588 178736 176594
rect 178684 176530 178736 176536
rect 184020 176588 184072 176594
rect 184020 176530 184072 176536
rect 193692 176526 193720 178092
rect 204916 176526 204944 200126
rect 212276 197962 212304 200330
rect 221372 200320 221424 200326
rect 221372 200262 221424 200268
rect 212060 197934 212304 197962
rect 221384 197962 221412 200262
rect 232596 200252 232648 200258
rect 232596 200194 232648 200200
rect 231032 200184 231084 200190
rect 231032 200126 231084 200132
rect 232504 200184 232556 200190
rect 232504 200126 232556 200132
rect 231044 197962 231072 200126
rect 221384 197934 221720 197962
rect 231044 197934 231380 197962
rect 209686 188320 209742 188329
rect 209686 188255 209742 188264
rect 205638 187640 205694 187649
rect 205638 187575 205694 187584
rect 205652 179314 205680 187575
rect 209700 179382 209728 188255
rect 209688 179376 209740 179382
rect 209688 179318 209740 179324
rect 205640 179308 205692 179314
rect 205640 179250 205692 179256
rect 231676 179308 231728 179314
rect 231676 179250 231728 179256
rect 231688 178786 231716 179250
rect 231380 178758 231716 178786
rect 211724 178078 212060 178106
rect 221720 178078 222056 178106
rect 211724 176594 211752 178078
rect 222028 176594 222056 178078
rect 232516 176594 232544 200126
rect 232608 179314 232636 200194
rect 232700 179926 232728 200330
rect 233238 187640 233294 187649
rect 233238 187575 233294 187584
rect 232688 179920 232740 179926
rect 232688 179862 232740 179868
rect 232596 179308 232648 179314
rect 232596 179250 232648 179256
rect 233252 179246 233280 187575
rect 233240 179240 233292 179246
rect 233240 179182 233292 179188
rect 211712 176588 211764 176594
rect 211712 176530 211764 176536
rect 222016 176588 222068 176594
rect 222016 176530 222068 176536
rect 232504 176588 232556 176594
rect 232504 176530 232556 176536
rect 81992 176520 82044 176526
rect 81992 176462 82044 176468
rect 94504 176520 94556 176526
rect 94504 176462 94556 176468
rect 109684 176520 109736 176526
rect 109684 176462 109736 176468
rect 120724 176520 120776 176526
rect 120724 176462 120776 176468
rect 137652 176520 137704 176526
rect 137652 176462 137704 176468
rect 148324 176520 148376 176526
rect 148324 176462 148376 176468
rect 193680 176520 193732 176526
rect 193680 176462 193732 176468
rect 204904 176520 204956 176526
rect 204904 176462 204956 176468
rect 212264 172780 212316 172786
rect 212264 172722 212316 172728
rect 232688 172780 232740 172786
rect 232688 172722 232740 172728
rect 148416 172712 148468 172718
rect 148416 172654 148468 172660
rect 165620 172712 165672 172718
rect 165620 172654 165672 172660
rect 175464 172712 175516 172718
rect 175464 172654 175516 172660
rect 193680 172712 193732 172718
rect 193680 172654 193732 172660
rect 203524 172712 203576 172718
rect 203524 172654 203576 172660
rect 81440 172644 81492 172650
rect 81440 172586 81492 172592
rect 91468 172644 91520 172650
rect 91468 172586 91520 172592
rect 109684 172644 109736 172650
rect 109684 172586 109736 172592
rect 119436 172644 119488 172650
rect 119436 172586 119488 172592
rect 137652 172644 137704 172650
rect 137652 172586 137704 172592
rect 81452 170898 81480 172586
rect 91100 172576 91152 172582
rect 91100 172518 91152 172524
rect 91112 170898 91140 172518
rect 81452 170870 81696 170898
rect 91112 170870 91356 170898
rect 71884 170326 72036 170354
rect 71044 148980 71096 148986
rect 71044 148922 71096 148928
rect 71884 148918 71912 170326
rect 91480 151722 91508 172586
rect 94504 172576 94556 172582
rect 94504 172518 94556 172524
rect 93858 160576 93914 160585
rect 93858 160511 93914 160520
rect 91356 151694 91508 151722
rect 93872 151706 93900 160511
rect 93860 151700 93912 151706
rect 93860 151642 93912 151648
rect 72036 151014 72096 151042
rect 81696 151014 82032 151042
rect 71872 148912 71924 148918
rect 71872 148854 71924 148860
rect 72068 148850 72096 151014
rect 82004 148850 82032 151014
rect 94516 148850 94544 172518
rect 109696 170884 109724 172586
rect 119344 172576 119396 172582
rect 119344 172518 119396 172524
rect 119356 170884 119384 172518
rect 99484 170326 100050 170354
rect 97906 161256 97962 161265
rect 97906 161191 97962 161200
rect 97920 151706 97948 161191
rect 97908 151700 97960 151706
rect 97908 151642 97960 151648
rect 99484 148850 99512 170326
rect 119448 151722 119476 172586
rect 120724 172576 120776 172582
rect 120724 172518 120776 172524
rect 119370 151694 119476 151722
rect 100036 148918 100064 151028
rect 100024 148912 100076 148918
rect 100024 148854 100076 148860
rect 109696 148850 109724 151028
rect 120736 148850 120764 172518
rect 137664 170884 137692 172586
rect 147312 172576 147364 172582
rect 147312 172518 147364 172524
rect 148324 172576 148376 172582
rect 148324 172518 148376 172524
rect 147324 170884 147352 172518
rect 127084 170326 128018 170354
rect 126886 161256 126942 161265
rect 126886 161191 126942 161200
rect 121458 160576 121514 160585
rect 121458 160511 121514 160520
rect 121472 151774 121500 160511
rect 126900 151774 126928 161191
rect 121460 151768 121512 151774
rect 121460 151710 121512 151716
rect 126888 151768 126940 151774
rect 126888 151710 126940 151716
rect 127084 148850 127112 170326
rect 147680 156664 147732 156670
rect 147680 156606 147732 156612
rect 147692 151722 147720 156606
rect 147338 151694 147720 151722
rect 128004 148918 128032 151028
rect 127992 148912 128044 148918
rect 127992 148854 128044 148860
rect 137664 148850 137692 151028
rect 148336 148850 148364 172518
rect 148428 156670 148456 172654
rect 156328 172644 156380 172650
rect 156328 172586 156380 172592
rect 156340 170898 156368 172586
rect 165632 171134 165660 172654
rect 175280 172576 175332 172582
rect 175280 172518 175332 172524
rect 175292 171134 175320 172518
rect 165632 171106 165706 171134
rect 175292 171106 175366 171134
rect 156032 170870 156368 170898
rect 165678 170884 165706 171106
rect 175338 170884 175366 171106
rect 154486 161256 154542 161265
rect 154486 161191 154542 161200
rect 149058 160576 149114 160585
rect 149058 160511 149114 160520
rect 148416 156664 148468 156670
rect 148416 156606 148468 156612
rect 149072 151706 149100 160511
rect 154500 151706 154528 161191
rect 175476 151722 175504 172654
rect 178684 172644 178736 172650
rect 178684 172586 178736 172592
rect 177304 172576 177356 172582
rect 177304 172518 177356 172524
rect 149060 151700 149112 151706
rect 149060 151642 149112 151648
rect 154488 151700 154540 151706
rect 175352 151694 175504 151722
rect 154488 151642 154540 151648
rect 156032 151014 156092 151042
rect 165692 151014 166028 151042
rect 156064 148918 156092 151014
rect 166000 148918 166028 151014
rect 177316 148918 177344 172518
rect 178038 160576 178094 160585
rect 178038 160511 178094 160520
rect 178052 151774 178080 160511
rect 178040 151768 178092 151774
rect 178040 151710 178092 151716
rect 178696 149054 178724 172586
rect 193692 170884 193720 172654
rect 203340 172576 203392 172582
rect 203340 172518 203392 172524
rect 203352 170884 203380 172518
rect 183664 170326 184046 170354
rect 182086 161256 182142 161265
rect 182086 161191 182142 161200
rect 182100 151638 182128 161191
rect 182088 151632 182140 151638
rect 182088 151574 182140 151580
rect 178684 149048 178736 149054
rect 178684 148990 178736 148996
rect 183664 148918 183692 170326
rect 203536 151722 203564 172654
rect 204904 172576 204956 172582
rect 204904 172518 204956 172524
rect 203366 151694 203564 151722
rect 184032 149054 184060 151028
rect 184020 149048 184072 149054
rect 184020 148990 184072 148996
rect 156052 148912 156104 148918
rect 156052 148854 156104 148860
rect 165988 148912 166040 148918
rect 165988 148854 166040 148860
rect 177304 148912 177356 148918
rect 177304 148854 177356 148860
rect 183652 148912 183704 148918
rect 183652 148854 183704 148860
rect 193692 148850 193720 151028
rect 204916 148850 204944 172518
rect 212276 170898 212304 172722
rect 221372 172712 221424 172718
rect 221372 172654 221424 172660
rect 212060 170870 212304 170898
rect 221384 170898 221412 172654
rect 232596 172644 232648 172650
rect 232596 172586 232648 172592
rect 231032 172576 231084 172582
rect 231032 172518 231084 172524
rect 232504 172576 232556 172582
rect 232504 172518 232556 172524
rect 231044 170898 231072 172518
rect 221384 170870 221720 170898
rect 231044 170870 231380 170898
rect 209686 161256 209742 161265
rect 209686 161191 209742 161200
rect 205638 160576 205694 160585
rect 205638 160511 205694 160520
rect 205652 151706 205680 160511
rect 209700 151774 209728 161191
rect 209688 151768 209740 151774
rect 209688 151710 209740 151716
rect 231380 151706 231716 151722
rect 205640 151700 205692 151706
rect 231380 151700 231728 151706
rect 231380 151694 231676 151700
rect 205640 151642 205692 151648
rect 231676 151642 231728 151648
rect 211724 151014 212060 151042
rect 221720 151014 222056 151042
rect 211724 148918 211752 151014
rect 222028 148918 222056 151014
rect 232516 148918 232544 172518
rect 232608 151706 232636 172586
rect 232700 152590 232728 172722
rect 233238 160576 233294 160585
rect 233238 160511 233294 160520
rect 232688 152584 232740 152590
rect 232688 152526 232740 152532
rect 232596 151700 232648 151706
rect 232596 151642 232648 151648
rect 233252 151638 233280 160511
rect 233240 151632 233292 151638
rect 233240 151574 233292 151580
rect 211712 148912 211764 148918
rect 211712 148854 211764 148860
rect 222016 148912 222068 148918
rect 222016 148854 222068 148860
rect 232504 148912 232556 148918
rect 232504 148854 232556 148860
rect 72056 148844 72108 148850
rect 72056 148786 72108 148792
rect 81992 148844 82044 148850
rect 81992 148786 82044 148792
rect 94504 148844 94556 148850
rect 94504 148786 94556 148792
rect 99472 148844 99524 148850
rect 99472 148786 99524 148792
rect 109684 148844 109736 148850
rect 109684 148786 109736 148792
rect 120724 148844 120776 148850
rect 120724 148786 120776 148792
rect 127072 148844 127124 148850
rect 127072 148786 127124 148792
rect 137652 148844 137704 148850
rect 137652 148786 137704 148792
rect 148324 148844 148376 148850
rect 148324 148786 148376 148792
rect 193680 148844 193732 148850
rect 193680 148786 193732 148792
rect 204904 148844 204956 148850
rect 204904 148786 204956 148792
rect 71044 146532 71096 146538
rect 71044 146474 71096 146480
rect 212356 146532 212408 146538
rect 212356 146474 212408 146480
rect 232688 146532 232740 146538
rect 232688 146474 232740 146480
rect 69664 146328 69716 146334
rect 69664 146270 69716 146276
rect 69676 122602 69704 146270
rect 70306 134328 70362 134337
rect 70306 134263 70362 134272
rect 70320 125594 70348 134263
rect 70308 125588 70360 125594
rect 70308 125530 70360 125536
rect 69664 122596 69716 122602
rect 69664 122538 69716 122544
rect 70306 107264 70362 107273
rect 70306 107199 70362 107208
rect 70320 97850 70348 107199
rect 70308 97844 70360 97850
rect 70308 97786 70360 97792
rect 71056 95130 71084 146474
rect 148416 146464 148468 146470
rect 148416 146406 148468 146412
rect 165712 146464 165764 146470
rect 165712 146406 165764 146412
rect 175464 146464 175516 146470
rect 175464 146406 175516 146412
rect 193680 146464 193732 146470
rect 193680 146406 193732 146412
rect 203524 146464 203576 146470
rect 203524 146406 203576 146412
rect 81440 146396 81492 146402
rect 81440 146338 81492 146344
rect 91468 146396 91520 146402
rect 91468 146338 91520 146344
rect 109684 146396 109736 146402
rect 109684 146338 109736 146344
rect 119436 146396 119488 146402
rect 119436 146338 119488 146344
rect 137652 146396 137704 146402
rect 137652 146338 137704 146344
rect 81452 143970 81480 146338
rect 91100 146328 91152 146334
rect 91100 146270 91152 146276
rect 91112 143970 91140 146270
rect 81452 143942 81696 143970
rect 91112 143942 91356 143970
rect 71884 143262 72036 143290
rect 71884 122670 71912 143262
rect 91480 124794 91508 146338
rect 94504 146328 94556 146334
rect 94504 146270 94556 146276
rect 93858 133648 93914 133657
rect 93858 133583 93914 133592
rect 93872 125526 93900 133583
rect 93860 125520 93912 125526
rect 93860 125462 93912 125468
rect 91356 124766 91508 124794
rect 72022 123842 72050 124100
rect 81696 124086 82032 124114
rect 71976 123814 72050 123842
rect 71872 122664 71924 122670
rect 71872 122606 71924 122612
rect 71976 122602 72004 123814
rect 82004 122602 82032 124086
rect 94516 122602 94544 146270
rect 109696 143956 109724 146338
rect 119344 146328 119396 146334
rect 119344 146270 119396 146276
rect 119356 143956 119384 146270
rect 99484 143262 100050 143290
rect 97906 134328 97962 134337
rect 97906 134263 97962 134272
rect 97920 125526 97948 134263
rect 97908 125520 97960 125526
rect 97908 125462 97960 125468
rect 99484 122602 99512 143262
rect 119448 124794 119476 146338
rect 120724 146328 120776 146334
rect 120724 146270 120776 146276
rect 119370 124766 119476 124794
rect 100036 122670 100064 124100
rect 100024 122664 100076 122670
rect 100024 122606 100076 122612
rect 109696 122602 109724 124100
rect 120736 122602 120764 146270
rect 137664 143956 137692 146338
rect 147312 146328 147364 146334
rect 147312 146270 147364 146276
rect 148324 146328 148376 146334
rect 148324 146270 148376 146276
rect 147324 143956 147352 146270
rect 127084 143262 128018 143290
rect 126886 134328 126942 134337
rect 126886 134263 126942 134272
rect 121458 133648 121514 133657
rect 121458 133583 121514 133592
rect 121472 125594 121500 133583
rect 126900 125594 126928 134263
rect 121460 125588 121512 125594
rect 121460 125530 121512 125536
rect 126888 125588 126940 125594
rect 126888 125530 126940 125536
rect 127084 122602 127112 143262
rect 147680 128308 147732 128314
rect 147680 128250 147732 128256
rect 147692 124794 147720 128250
rect 147338 124766 147720 124794
rect 128004 122670 128032 124100
rect 127992 122664 128044 122670
rect 127992 122606 128044 122612
rect 137664 122602 137692 124100
rect 148336 122602 148364 146270
rect 148428 128314 148456 146406
rect 156328 146396 156380 146402
rect 156328 146338 156380 146344
rect 156340 143970 156368 146338
rect 156032 143942 156368 143970
rect 165724 143834 165752 146406
rect 175372 146328 175424 146334
rect 175372 146270 175424 146276
rect 175384 143834 175412 146270
rect 165692 143806 165752 143834
rect 175352 143806 175412 143834
rect 154486 134328 154542 134337
rect 154486 134263 154542 134272
rect 149058 133648 149114 133657
rect 149058 133583 149114 133592
rect 148416 128308 148468 128314
rect 148416 128250 148468 128256
rect 149072 125526 149100 133583
rect 154500 125526 154528 134263
rect 149060 125520 149112 125526
rect 149060 125462 149112 125468
rect 154488 125520 154540 125526
rect 154488 125462 154540 125468
rect 175476 124794 175504 146406
rect 178684 146396 178736 146402
rect 178684 146338 178736 146344
rect 177304 146328 177356 146334
rect 177304 146270 177356 146276
rect 175352 124766 175504 124794
rect 156018 123842 156046 124100
rect 165692 124086 166028 124114
rect 155972 123814 156046 123842
rect 155972 122670 156000 123814
rect 166000 122670 166028 124086
rect 177316 122670 177344 146270
rect 178038 133648 178094 133657
rect 178038 133583 178094 133592
rect 178052 125594 178080 133583
rect 178040 125588 178092 125594
rect 178040 125530 178092 125536
rect 178696 122806 178724 146338
rect 193692 143956 193720 146406
rect 203340 146328 203392 146334
rect 203340 146270 203392 146276
rect 203352 143956 203380 146270
rect 183664 143262 184046 143290
rect 182086 134328 182142 134337
rect 182086 134263 182142 134272
rect 182100 125458 182128 134263
rect 182088 125452 182140 125458
rect 182088 125394 182140 125400
rect 178684 122800 178736 122806
rect 178684 122742 178736 122748
rect 183664 122670 183692 143262
rect 203536 124794 203564 146406
rect 204904 146328 204956 146334
rect 204904 146270 204956 146276
rect 203366 124766 203564 124794
rect 184032 122806 184060 124100
rect 184020 122800 184072 122806
rect 184020 122742 184072 122748
rect 155960 122664 156012 122670
rect 155960 122606 156012 122612
rect 165988 122664 166040 122670
rect 165988 122606 166040 122612
rect 177304 122664 177356 122670
rect 177304 122606 177356 122612
rect 183652 122664 183704 122670
rect 183652 122606 183704 122612
rect 193692 122602 193720 124100
rect 204916 122602 204944 146270
rect 212368 143970 212396 146474
rect 221372 146464 221424 146470
rect 221372 146406 221424 146412
rect 212060 143942 212396 143970
rect 221384 143970 221412 146406
rect 232504 146396 232556 146402
rect 232504 146338 232556 146344
rect 231032 146328 231084 146334
rect 231032 146270 231084 146276
rect 231044 143970 231072 146270
rect 221384 143942 221720 143970
rect 231044 143942 231380 143970
rect 209686 134328 209742 134337
rect 209686 134263 209742 134272
rect 205638 133648 205694 133657
rect 205638 133583 205694 133592
rect 205652 125526 205680 133583
rect 209700 125594 209728 134263
rect 209688 125588 209740 125594
rect 209688 125530 209740 125536
rect 205640 125520 205692 125526
rect 205640 125462 205692 125468
rect 211724 124086 212060 124114
rect 221720 124086 221964 124114
rect 231380 124086 231624 124114
rect 211724 122670 211752 124086
rect 221936 122670 221964 124086
rect 231596 122806 231624 124086
rect 232516 122806 232544 146338
rect 232596 146328 232648 146334
rect 232596 146270 232648 146276
rect 231584 122800 231636 122806
rect 231584 122742 231636 122748
rect 232504 122800 232556 122806
rect 232504 122742 232556 122748
rect 232608 122670 232636 146270
rect 232700 126954 232728 146474
rect 233238 133648 233294 133657
rect 233238 133583 233294 133592
rect 232688 126948 232740 126954
rect 232688 126890 232740 126896
rect 233252 125458 233280 133583
rect 233240 125452 233292 125458
rect 233240 125394 233292 125400
rect 211712 122664 211764 122670
rect 211712 122606 211764 122612
rect 221924 122664 221976 122670
rect 221924 122606 221976 122612
rect 232596 122664 232648 122670
rect 232596 122606 232648 122612
rect 71964 122596 72016 122602
rect 71964 122538 72016 122544
rect 81992 122596 82044 122602
rect 81992 122538 82044 122544
rect 94504 122596 94556 122602
rect 94504 122538 94556 122544
rect 99472 122596 99524 122602
rect 99472 122538 99524 122544
rect 109684 122596 109736 122602
rect 109684 122538 109736 122544
rect 120724 122596 120776 122602
rect 120724 122538 120776 122544
rect 127072 122596 127124 122602
rect 127072 122538 127124 122544
rect 137652 122596 137704 122602
rect 137652 122538 137704 122544
rect 148324 122596 148376 122602
rect 148324 122538 148376 122544
rect 193680 122596 193732 122602
rect 193680 122538 193732 122544
rect 204904 122596 204956 122602
rect 204904 122538 204956 122544
rect 148324 118924 148376 118930
rect 148324 118866 148376 118872
rect 165712 118924 165764 118930
rect 165712 118866 165764 118872
rect 175464 118924 175516 118930
rect 175464 118866 175516 118872
rect 193680 118924 193732 118930
rect 193680 118866 193732 118872
rect 203524 118924 203576 118930
rect 203524 118866 203576 118872
rect 221372 118924 221424 118930
rect 221372 118866 221424 118872
rect 81440 118856 81492 118862
rect 81440 118798 81492 118804
rect 91468 118856 91520 118862
rect 91468 118798 91520 118804
rect 109684 118856 109736 118862
rect 109684 118798 109736 118804
rect 119436 118856 119488 118862
rect 119436 118798 119488 118804
rect 137652 118856 137704 118862
rect 137652 118798 137704 118804
rect 81452 116906 81480 118798
rect 91100 118788 91152 118794
rect 91100 118730 91152 118736
rect 91112 116906 91140 118730
rect 81452 116878 81696 116906
rect 91112 116878 91356 116906
rect 71884 116334 72036 116362
rect 71044 95124 71096 95130
rect 71044 95066 71096 95072
rect 71884 95062 71912 116334
rect 91480 97730 91508 118798
rect 94504 118788 94556 118794
rect 94504 118730 94556 118736
rect 93858 106584 93914 106593
rect 93858 106519 93914 106528
rect 93872 97918 93900 106519
rect 93860 97912 93912 97918
rect 93860 97854 93912 97860
rect 91356 97702 91508 97730
rect 72036 97022 72096 97050
rect 81696 97022 82032 97050
rect 71872 95056 71924 95062
rect 71872 94998 71924 95004
rect 72068 94994 72096 97022
rect 82004 94994 82032 97022
rect 94516 94994 94544 118730
rect 109696 116892 109724 118798
rect 119344 118788 119396 118794
rect 119344 118730 119396 118736
rect 119356 116892 119384 118730
rect 99484 116334 100050 116362
rect 97906 107264 97962 107273
rect 97906 107199 97962 107208
rect 97920 97986 97948 107199
rect 97908 97980 97960 97986
rect 97908 97922 97960 97928
rect 99484 94994 99512 116334
rect 119448 97730 119476 118798
rect 120724 118788 120776 118794
rect 120724 118730 120776 118736
rect 119370 97702 119476 97730
rect 100036 95062 100064 97036
rect 100024 95056 100076 95062
rect 100024 94998 100076 95004
rect 109696 94994 109724 97036
rect 120736 94994 120764 118730
rect 137664 116892 137692 118798
rect 147312 118788 147364 118794
rect 147312 118730 147364 118736
rect 147324 116892 147352 118730
rect 127084 116334 128018 116362
rect 126886 107264 126942 107273
rect 126886 107199 126942 107208
rect 121458 106584 121514 106593
rect 121458 106519 121514 106528
rect 121472 97850 121500 106519
rect 126900 97918 126928 107199
rect 126888 97912 126940 97918
rect 126888 97854 126940 97860
rect 121460 97844 121512 97850
rect 121460 97786 121512 97792
rect 127084 94994 127112 116334
rect 148336 103514 148364 118866
rect 156328 118856 156380 118862
rect 156328 118798 156380 118804
rect 148416 118788 148468 118794
rect 148416 118730 148468 118736
rect 147784 103486 148364 103514
rect 147784 97730 147812 103486
rect 147338 97702 147812 97730
rect 128004 95062 128032 97036
rect 127992 95056 128044 95062
rect 127992 94998 128044 95004
rect 137664 94994 137692 97036
rect 148428 94994 148456 118730
rect 156340 116906 156368 118798
rect 156032 116878 156368 116906
rect 165724 116770 165752 118866
rect 175372 118788 175424 118794
rect 175372 118730 175424 118736
rect 175384 116770 175412 118730
rect 165692 116742 165752 116770
rect 175352 116742 175412 116770
rect 154486 107264 154542 107273
rect 154486 107199 154542 107208
rect 149058 106584 149114 106593
rect 149058 106519 149114 106528
rect 149072 97986 149100 106519
rect 154500 97986 154528 107199
rect 149060 97980 149112 97986
rect 149060 97922 149112 97928
rect 154488 97980 154540 97986
rect 154488 97922 154540 97928
rect 175476 97730 175504 118866
rect 178684 118856 178736 118862
rect 178684 118798 178736 118804
rect 177304 118788 177356 118794
rect 177304 118730 177356 118736
rect 175352 97702 175504 97730
rect 156032 97022 156092 97050
rect 165692 97022 166028 97050
rect 156064 95062 156092 97022
rect 166000 95062 166028 97022
rect 177316 95062 177344 118730
rect 178038 106584 178094 106593
rect 178038 106519 178094 106528
rect 178052 97918 178080 106519
rect 178040 97912 178092 97918
rect 178040 97854 178092 97860
rect 178696 95198 178724 118798
rect 193692 116892 193720 118866
rect 203340 118788 203392 118794
rect 203340 118730 203392 118736
rect 203352 116892 203380 118730
rect 183664 116334 184046 116362
rect 182086 107264 182142 107273
rect 182086 107199 182142 107208
rect 182100 97918 182128 107199
rect 182088 97912 182140 97918
rect 182088 97854 182140 97860
rect 178684 95192 178736 95198
rect 178684 95134 178736 95140
rect 183664 95062 183692 116334
rect 203536 97730 203564 118866
rect 204904 118788 204956 118794
rect 204904 118730 204956 118736
rect 203366 97702 203564 97730
rect 184032 95198 184060 97036
rect 184020 95192 184072 95198
rect 184020 95134 184072 95140
rect 156052 95056 156104 95062
rect 156052 94998 156104 95004
rect 165988 95056 166040 95062
rect 165988 94998 166040 95004
rect 177304 95056 177356 95062
rect 177304 94998 177356 95004
rect 183652 95056 183704 95062
rect 183652 94998 183704 95004
rect 193692 94994 193720 97036
rect 204916 94994 204944 118730
rect 212356 118720 212408 118726
rect 212356 118662 212408 118668
rect 212368 116906 212396 118662
rect 212060 116878 212396 116906
rect 221384 116906 221412 118866
rect 232596 118856 232648 118862
rect 232596 118798 232648 118804
rect 231032 118788 231084 118794
rect 231032 118730 231084 118736
rect 232504 118788 232556 118794
rect 232504 118730 232556 118736
rect 231044 116906 231072 118730
rect 221384 116878 221720 116906
rect 231044 116878 231380 116906
rect 209686 107264 209742 107273
rect 209686 107199 209742 107208
rect 205638 106584 205694 106593
rect 205638 106519 205694 106528
rect 205652 97986 205680 106519
rect 209700 97986 209728 107199
rect 205640 97980 205692 97986
rect 205640 97922 205692 97928
rect 209688 97980 209740 97986
rect 209688 97922 209740 97928
rect 231676 97844 231728 97850
rect 231676 97786 231728 97792
rect 231688 97730 231716 97786
rect 231380 97702 231716 97730
rect 211724 97022 212060 97050
rect 221720 97022 222056 97050
rect 211724 95062 211752 97022
rect 222028 95062 222056 97022
rect 232516 95062 232544 118730
rect 232608 97850 232636 118798
rect 232688 118720 232740 118726
rect 232688 118662 232740 118668
rect 232700 98258 232728 118662
rect 233238 106584 233294 106593
rect 233238 106519 233294 106528
rect 232688 98252 232740 98258
rect 232688 98194 232740 98200
rect 233252 97918 233280 106519
rect 233240 97912 233292 97918
rect 233240 97854 233292 97860
rect 232596 97844 232648 97850
rect 232596 97786 232648 97792
rect 211712 95056 211764 95062
rect 211712 94998 211764 95004
rect 222016 95056 222068 95062
rect 222016 94998 222068 95004
rect 232504 95056 232556 95062
rect 232504 94998 232556 95004
rect 72056 94988 72108 94994
rect 72056 94930 72108 94936
rect 81992 94988 82044 94994
rect 81992 94930 82044 94936
rect 94504 94988 94556 94994
rect 94504 94930 94556 94936
rect 99472 94988 99524 94994
rect 99472 94930 99524 94936
rect 109684 94988 109736 94994
rect 109684 94930 109736 94936
rect 120724 94988 120776 94994
rect 120724 94930 120776 94936
rect 127072 94988 127124 94994
rect 127072 94930 127124 94936
rect 137652 94988 137704 94994
rect 137652 94930 137704 94936
rect 148416 94988 148468 94994
rect 148416 94930 148468 94936
rect 193680 94988 193732 94994
rect 193680 94930 193732 94936
rect 204904 94988 204956 94994
rect 204904 94930 204956 94936
rect 71044 91316 71096 91322
rect 71044 91258 71096 91264
rect 212356 91316 212408 91322
rect 212356 91258 212408 91264
rect 232688 91316 232740 91322
rect 232688 91258 232740 91264
rect 69664 91112 69716 91118
rect 69664 91054 69716 91060
rect 69676 68882 69704 91054
rect 70308 88392 70360 88398
rect 70308 88334 70360 88340
rect 70320 80345 70348 88334
rect 70306 80336 70362 80345
rect 70306 80271 70362 80280
rect 69664 68876 69716 68882
rect 69664 68818 69716 68824
rect 70306 53272 70362 53281
rect 70306 53207 70362 53216
rect 70320 44130 70348 53207
rect 70308 44124 70360 44130
rect 70308 44066 70360 44072
rect 71056 41342 71084 91258
rect 148324 91248 148376 91254
rect 148324 91190 148376 91196
rect 165712 91248 165764 91254
rect 165712 91190 165764 91196
rect 175464 91248 175516 91254
rect 175464 91190 175516 91196
rect 193680 91248 193732 91254
rect 193680 91190 193732 91196
rect 203524 91248 203576 91254
rect 203524 91190 203576 91196
rect 81440 91180 81492 91186
rect 81440 91122 81492 91128
rect 91468 91180 91520 91186
rect 91468 91122 91520 91128
rect 109684 91180 109736 91186
rect 109684 91122 109736 91128
rect 119436 91180 119488 91186
rect 119436 91122 119488 91128
rect 137652 91180 137704 91186
rect 137652 91122 137704 91128
rect 81452 89978 81480 91122
rect 91100 91112 91152 91118
rect 91100 91054 91152 91060
rect 91112 89978 91140 91054
rect 81452 89950 81696 89978
rect 91112 89950 91356 89978
rect 71884 89270 72036 89298
rect 71884 68950 71912 89270
rect 91480 70666 91508 91122
rect 94504 91112 94556 91118
rect 94504 91054 94556 91060
rect 93860 88460 93912 88466
rect 93860 88402 93912 88408
rect 93872 79665 93900 88402
rect 93858 79656 93914 79665
rect 93858 79591 93914 79600
rect 91356 70638 91508 70666
rect 72036 70094 72096 70122
rect 81696 70094 82032 70122
rect 72068 69018 72096 70094
rect 72056 69012 72108 69018
rect 72056 68954 72108 68960
rect 71872 68944 71924 68950
rect 71872 68886 71924 68892
rect 82004 68882 82032 70094
rect 94516 68882 94544 91054
rect 109696 89964 109724 91122
rect 119344 91112 119396 91118
rect 119344 91054 119396 91060
rect 119356 89964 119384 91054
rect 99484 89270 100050 89298
rect 97906 80336 97962 80345
rect 97906 80271 97962 80280
rect 97920 71738 97948 80271
rect 97908 71732 97960 71738
rect 97908 71674 97960 71680
rect 99484 69018 99512 89270
rect 119448 70666 119476 91122
rect 120724 91112 120776 91118
rect 120724 91054 120776 91060
rect 119370 70638 119476 70666
rect 99472 69012 99524 69018
rect 99472 68954 99524 68960
rect 100036 68950 100064 70108
rect 100024 68944 100076 68950
rect 100024 68886 100076 68892
rect 109696 68882 109724 70108
rect 120736 68882 120764 91054
rect 137664 89964 137692 91122
rect 147312 91112 147364 91118
rect 147312 91054 147364 91060
rect 147324 89964 147352 91054
rect 127084 89270 128018 89298
rect 121460 88392 121512 88398
rect 121460 88334 121512 88340
rect 126888 88392 126940 88398
rect 126888 88334 126940 88340
rect 121472 79665 121500 88334
rect 126900 80345 126928 88334
rect 126886 80336 126942 80345
rect 126886 80271 126942 80280
rect 121458 79656 121514 79665
rect 121458 79591 121514 79600
rect 127084 69018 127112 89270
rect 148336 74534 148364 91190
rect 156328 91180 156380 91186
rect 156328 91122 156380 91128
rect 148416 91112 148468 91118
rect 148416 91054 148468 91060
rect 147784 74506 148364 74534
rect 147784 70666 147812 74506
rect 147338 70638 147812 70666
rect 127072 69012 127124 69018
rect 127072 68954 127124 68960
rect 128004 68950 128032 70108
rect 127992 68944 128044 68950
rect 127992 68886 128044 68892
rect 137664 68882 137692 70108
rect 148428 68882 148456 91054
rect 156340 89978 156368 91122
rect 156032 89950 156368 89978
rect 165724 89842 165752 91190
rect 175372 91112 175424 91118
rect 175372 91054 175424 91060
rect 175384 89842 175412 91054
rect 165692 89814 165752 89842
rect 175352 89814 175412 89842
rect 154488 88460 154540 88466
rect 154488 88402 154540 88408
rect 154500 80345 154528 88402
rect 154486 80336 154542 80345
rect 154486 80271 154542 80280
rect 149058 79656 149114 79665
rect 149058 79591 149114 79600
rect 149072 71738 149100 79591
rect 149060 71732 149112 71738
rect 149060 71674 149112 71680
rect 175476 70666 175504 91190
rect 178684 91180 178736 91186
rect 178684 91122 178736 91128
rect 177304 91112 177356 91118
rect 177304 91054 177356 91060
rect 175352 70638 175504 70666
rect 156032 70094 156092 70122
rect 165692 70094 166028 70122
rect 156064 68950 156092 70094
rect 166000 68950 166028 70094
rect 177316 68950 177344 91054
rect 178040 88392 178092 88398
rect 178040 88334 178092 88340
rect 178052 79665 178080 88334
rect 178038 79656 178094 79665
rect 178038 79591 178094 79600
rect 178696 68950 178724 91122
rect 193692 89964 193720 91190
rect 203340 91112 203392 91118
rect 203340 91054 203392 91060
rect 203352 89964 203380 91054
rect 183664 89270 184046 89298
rect 182086 80336 182142 80345
rect 182086 80271 182142 80280
rect 182100 71738 182128 80271
rect 182088 71732 182140 71738
rect 182088 71674 182140 71680
rect 183664 69018 183692 89270
rect 203536 70666 203564 91190
rect 204904 91112 204956 91118
rect 204904 91054 204956 91060
rect 203366 70638 203564 70666
rect 183652 69012 183704 69018
rect 183652 68954 183704 68960
rect 184032 68950 184060 70108
rect 156052 68944 156104 68950
rect 156052 68886 156104 68892
rect 165988 68944 166040 68950
rect 165988 68886 166040 68892
rect 177304 68944 177356 68950
rect 177304 68886 177356 68892
rect 178684 68944 178736 68950
rect 178684 68886 178736 68892
rect 184020 68944 184072 68950
rect 184020 68886 184072 68892
rect 193692 68882 193720 70108
rect 204916 68882 204944 91054
rect 212368 89978 212396 91258
rect 221372 91248 221424 91254
rect 221372 91190 221424 91196
rect 212060 89950 212396 89978
rect 221384 89978 221412 91190
rect 232596 91180 232648 91186
rect 232596 91122 232648 91128
rect 231032 91112 231084 91118
rect 231032 91054 231084 91060
rect 232504 91112 232556 91118
rect 232504 91054 232556 91060
rect 231044 89978 231072 91054
rect 221384 89950 221720 89978
rect 231044 89950 231380 89978
rect 205640 88460 205692 88466
rect 205640 88402 205692 88408
rect 205652 79665 205680 88402
rect 209688 88392 209740 88398
rect 209688 88334 209740 88340
rect 209700 80345 209728 88334
rect 209686 80336 209742 80345
rect 209686 80271 209742 80280
rect 205638 79656 205694 79665
rect 205638 79591 205694 79600
rect 231676 71664 231728 71670
rect 231676 71606 231728 71612
rect 231688 70666 231716 71606
rect 231380 70638 231716 70666
rect 211724 70094 212060 70122
rect 221720 70094 222056 70122
rect 211724 68950 211752 70094
rect 222028 68950 222056 70094
rect 232516 68950 232544 91054
rect 232608 71670 232636 91122
rect 232700 72350 232728 91258
rect 233238 79656 233294 79665
rect 233238 79591 233294 79600
rect 232688 72344 232740 72350
rect 232688 72286 232740 72292
rect 233252 71738 233280 79591
rect 233240 71732 233292 71738
rect 233240 71674 233292 71680
rect 232596 71664 232648 71670
rect 232596 71606 232648 71612
rect 211712 68944 211764 68950
rect 211712 68886 211764 68892
rect 222016 68944 222068 68950
rect 222016 68886 222068 68892
rect 232504 68944 232556 68950
rect 232504 68886 232556 68892
rect 81992 68876 82044 68882
rect 81992 68818 82044 68824
rect 94504 68876 94556 68882
rect 94504 68818 94556 68824
rect 109684 68876 109736 68882
rect 109684 68818 109736 68824
rect 120724 68876 120776 68882
rect 120724 68818 120776 68824
rect 137652 68876 137704 68882
rect 137652 68818 137704 68824
rect 148416 68876 148468 68882
rect 148416 68818 148468 68824
rect 193680 68876 193732 68882
rect 193680 68818 193732 68824
rect 204904 68876 204956 68882
rect 204904 68818 204956 68824
rect 148416 65136 148468 65142
rect 148416 65078 148468 65084
rect 165620 65136 165672 65142
rect 165620 65078 165672 65084
rect 175464 65136 175516 65142
rect 175464 65078 175516 65084
rect 193680 65136 193732 65142
rect 193680 65078 193732 65084
rect 203524 65136 203576 65142
rect 203524 65078 203576 65084
rect 221372 65136 221424 65142
rect 221372 65078 221424 65084
rect 81440 65068 81492 65074
rect 81440 65010 81492 65016
rect 91468 65068 91520 65074
rect 91468 65010 91520 65016
rect 109684 65068 109736 65074
rect 109684 65010 109736 65016
rect 119436 65068 119488 65074
rect 119436 65010 119488 65016
rect 137652 65068 137704 65074
rect 137652 65010 137704 65016
rect 81452 62914 81480 65010
rect 91100 65000 91152 65006
rect 91100 64942 91152 64948
rect 91112 62914 91140 64942
rect 81452 62886 81696 62914
rect 91112 62886 91356 62914
rect 71884 62206 72036 62234
rect 71044 41336 71096 41342
rect 71044 41278 71096 41284
rect 71884 41274 71912 62206
rect 91480 43738 91508 65010
rect 94504 65000 94556 65006
rect 94504 64942 94556 64948
rect 93860 62144 93912 62150
rect 93860 62086 93912 62092
rect 93872 52601 93900 62086
rect 93858 52592 93914 52601
rect 93858 52527 93914 52536
rect 91356 43710 91508 43738
rect 72036 43030 72096 43058
rect 81696 43030 82032 43058
rect 71872 41268 71924 41274
rect 71872 41210 71924 41216
rect 72068 41206 72096 43030
rect 82004 41206 82032 43030
rect 94516 41206 94544 64942
rect 109696 62900 109724 65010
rect 119344 65000 119396 65006
rect 119344 64942 119396 64948
rect 119356 62900 119384 64942
rect 99484 62206 100050 62234
rect 97908 62144 97960 62150
rect 97908 62086 97960 62092
rect 97920 53281 97948 62086
rect 97906 53272 97962 53281
rect 97906 53207 97962 53216
rect 99484 41206 99512 62206
rect 119448 43738 119476 65010
rect 120724 65000 120776 65006
rect 120724 64942 120776 64948
rect 119370 43710 119476 43738
rect 100036 41274 100064 43044
rect 100024 41268 100076 41274
rect 100024 41210 100076 41216
rect 109696 41206 109724 43044
rect 120736 41206 120764 64942
rect 137664 62900 137692 65010
rect 147312 65000 147364 65006
rect 147312 64942 147364 64948
rect 148324 65000 148376 65006
rect 148324 64942 148376 64948
rect 147324 62900 147352 64942
rect 127084 62206 128018 62234
rect 126886 53272 126942 53281
rect 126886 53207 126942 53216
rect 121458 52592 121514 52601
rect 121458 52527 121514 52536
rect 121472 44130 121500 52527
rect 126900 44130 126928 53207
rect 121460 44124 121512 44130
rect 121460 44066 121512 44072
rect 126888 44124 126940 44130
rect 126888 44066 126940 44072
rect 127084 41206 127112 62206
rect 147680 50380 147732 50386
rect 147680 50322 147732 50328
rect 147692 43738 147720 50322
rect 147338 43710 147720 43738
rect 128004 41274 128032 43044
rect 127992 41268 128044 41274
rect 127992 41210 128044 41216
rect 137664 41206 137692 43044
rect 148336 41206 148364 64942
rect 148428 50386 148456 65078
rect 156328 65068 156380 65074
rect 156328 65010 156380 65016
rect 156340 62914 156368 65010
rect 165632 63186 165660 65078
rect 175280 65000 175332 65006
rect 175280 64942 175332 64948
rect 175292 63186 175320 64942
rect 165632 63158 165706 63186
rect 175292 63158 175366 63186
rect 156032 62886 156368 62914
rect 165678 62900 165706 63158
rect 175338 62900 175366 63158
rect 149060 62144 149112 62150
rect 149060 62086 149112 62092
rect 154488 62144 154540 62150
rect 154488 62086 154540 62092
rect 149072 52601 149100 62086
rect 154500 53281 154528 62086
rect 154486 53272 154542 53281
rect 154486 53207 154542 53216
rect 149058 52592 149114 52601
rect 149058 52527 149114 52536
rect 148416 50380 148468 50386
rect 148416 50322 148468 50328
rect 175476 43738 175504 65078
rect 178684 65068 178736 65074
rect 178684 65010 178736 65016
rect 177304 65000 177356 65006
rect 177304 64942 177356 64948
rect 175352 43710 175504 43738
rect 156032 43030 156092 43058
rect 165692 43030 166028 43058
rect 156064 41274 156092 43030
rect 166000 41274 166028 43030
rect 177316 41274 177344 64942
rect 178038 52592 178094 52601
rect 178038 52527 178094 52536
rect 178052 44130 178080 52527
rect 178040 44124 178092 44130
rect 178040 44066 178092 44072
rect 178696 41410 178724 65010
rect 193692 62900 193720 65078
rect 203340 65000 203392 65006
rect 203340 64942 203392 64948
rect 203352 62900 203380 64942
rect 182088 62212 182140 62218
rect 182088 62154 182140 62160
rect 183664 62206 184046 62234
rect 182100 53281 182128 62154
rect 182086 53272 182142 53281
rect 182086 53207 182142 53216
rect 178684 41404 178736 41410
rect 178684 41346 178736 41352
rect 183664 41274 183692 62206
rect 203536 43738 203564 65078
rect 204904 65000 204956 65006
rect 204904 64942 204956 64948
rect 203366 43710 203564 43738
rect 184032 41410 184060 43044
rect 184020 41404 184072 41410
rect 184020 41346 184072 41352
rect 156052 41268 156104 41274
rect 156052 41210 156104 41216
rect 165988 41268 166040 41274
rect 165988 41210 166040 41216
rect 177304 41268 177356 41274
rect 177304 41210 177356 41216
rect 183652 41268 183704 41274
rect 183652 41210 183704 41216
rect 193692 41206 193720 43044
rect 204916 41206 204944 64942
rect 212264 64932 212316 64938
rect 212264 64874 212316 64880
rect 212276 62914 212304 64874
rect 212060 62886 212304 62914
rect 221384 62914 221412 65078
rect 232504 65068 232556 65074
rect 232504 65010 232556 65016
rect 231032 65000 231084 65006
rect 231032 64942 231084 64948
rect 231044 62914 231072 64942
rect 221384 62886 221720 62914
rect 231044 62886 231380 62914
rect 205640 62144 205692 62150
rect 205640 62086 205692 62092
rect 205652 52601 205680 62086
rect 209686 53272 209742 53281
rect 209686 53207 209742 53216
rect 205638 52592 205694 52601
rect 205638 52527 205694 52536
rect 209700 44130 209728 53207
rect 232516 45554 232544 65010
rect 232596 65000 232648 65006
rect 232596 64942 232648 64948
rect 231872 45526 232544 45554
rect 209688 44124 209740 44130
rect 209688 44066 209740 44072
rect 231872 43874 231900 45526
rect 231780 43846 231900 43874
rect 231780 43738 231808 43846
rect 231380 43710 231808 43738
rect 211724 43030 212060 43058
rect 221720 43030 222056 43058
rect 211724 41274 211752 43030
rect 222028 41274 222056 43030
rect 232608 41274 232636 64942
rect 232688 64932 232740 64938
rect 232688 64874 232740 64880
rect 232700 44946 232728 64874
rect 233240 62212 233292 62218
rect 233240 62154 233292 62160
rect 233252 52601 233280 62154
rect 233238 52592 233294 52601
rect 233238 52527 233294 52536
rect 232688 44940 232740 44946
rect 232688 44882 232740 44888
rect 211712 41268 211764 41274
rect 211712 41210 211764 41216
rect 222016 41268 222068 41274
rect 222016 41210 222068 41216
rect 232596 41268 232648 41274
rect 232596 41210 232648 41216
rect 72056 41200 72108 41206
rect 72056 41142 72108 41148
rect 81992 41200 82044 41206
rect 81992 41142 82044 41148
rect 94504 41200 94556 41206
rect 94504 41142 94556 41148
rect 99472 41200 99524 41206
rect 99472 41142 99524 41148
rect 109684 41200 109736 41206
rect 109684 41142 109736 41148
rect 120724 41200 120776 41206
rect 120724 41142 120776 41148
rect 127072 41200 127124 41206
rect 127072 41142 127124 41148
rect 137652 41200 137704 41206
rect 137652 41142 137704 41148
rect 148324 41200 148376 41206
rect 148324 41142 148376 41148
rect 193680 41200 193732 41206
rect 193680 41142 193732 41148
rect 204904 41200 204956 41206
rect 204904 41142 204956 41148
rect 234632 38078 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 300136 700534 300164 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 429856 700398 429884 703520
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 494808 699718 494836 703520
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 490564 699712 490616 699718
rect 490564 699654 490616 699660
rect 494796 699712 494848 699718
rect 494796 699654 494848 699660
rect 296352 686112 296404 686118
rect 296352 686054 296404 686060
rect 316776 686112 316828 686118
rect 316776 686054 316828 686060
rect 408040 686112 408092 686118
rect 408040 686054 408092 686060
rect 428648 686112 428700 686118
rect 428648 686054 428700 686060
rect 260196 686044 260248 686050
rect 260196 685986 260248 685992
rect 277676 686044 277728 686050
rect 277676 685986 277728 685992
rect 287520 686044 287572 686050
rect 287520 685986 287572 685992
rect 249708 685976 249760 685982
rect 249708 685918 249760 685924
rect 249720 683876 249748 685918
rect 259368 685908 259420 685914
rect 259368 685850 259420 685856
rect 260104 685908 260156 685914
rect 260104 685850 260156 685856
rect 259380 683876 259408 685850
rect 238864 683318 240074 683346
rect 238668 683188 238720 683194
rect 238668 683130 238720 683136
rect 238680 674257 238708 683130
rect 238666 674248 238722 674257
rect 238666 674183 238722 674192
rect 238864 662250 238892 683318
rect 259736 668772 259788 668778
rect 259736 668714 259788 668720
rect 239772 665304 239824 665310
rect 239772 665246 239824 665252
rect 239784 664714 239812 665246
rect 259748 664714 259776 668714
rect 239784 664686 240074 664714
rect 259394 664686 259776 664714
rect 249536 664142 249734 664170
rect 249536 663794 249564 664142
rect 249536 663766 249656 663794
rect 249628 662318 249656 663766
rect 260116 662318 260144 685850
rect 260208 668778 260236 685986
rect 268016 685976 268068 685982
rect 268016 685918 268068 685924
rect 268028 683876 268056 685918
rect 277688 683876 277716 685986
rect 287336 685908 287388 685914
rect 287336 685850 287388 685856
rect 287348 683876 287376 685850
rect 266266 674248 266322 674257
rect 266266 674183 266322 674192
rect 262218 673568 262274 673577
rect 262218 673503 262274 673512
rect 260196 668772 260248 668778
rect 260196 668714 260248 668720
rect 262232 665174 262260 673503
rect 266280 665174 266308 674183
rect 262220 665168 262272 665174
rect 262220 665110 262272 665116
rect 266268 665168 266320 665174
rect 266268 665110 266320 665116
rect 287532 664714 287560 685986
rect 287704 685976 287756 685982
rect 287704 685918 287756 685924
rect 287716 665514 287744 685918
rect 289084 685908 289136 685914
rect 289084 685850 289136 685856
rect 287704 665508 287756 665514
rect 287704 665450 287756 665456
rect 287362 664686 287560 664714
rect 249616 662312 249668 662318
rect 249616 662254 249668 662260
rect 260104 662312 260156 662318
rect 260104 662254 260156 662260
rect 268028 662250 268056 664020
rect 277688 662386 277716 664020
rect 289096 662386 289124 685850
rect 296364 683890 296392 686054
rect 305368 686044 305420 686050
rect 305368 685986 305420 685992
rect 296056 683862 296392 683890
rect 305380 683890 305408 685986
rect 315488 685976 315540 685982
rect 315488 685918 315540 685924
rect 315028 685908 315080 685914
rect 315028 685850 315080 685856
rect 315040 683890 315068 685850
rect 305380 683862 305716 683890
rect 315040 683862 315376 683890
rect 289820 683188 289872 683194
rect 289820 683130 289872 683136
rect 293868 683188 293920 683194
rect 293868 683130 293920 683136
rect 289832 673577 289860 683130
rect 293880 674257 293908 683130
rect 293866 674248 293922 674257
rect 293866 674183 293922 674192
rect 289818 673568 289874 673577
rect 289818 673503 289874 673512
rect 295708 665508 295760 665514
rect 295708 665450 295760 665456
rect 295720 664714 295748 665450
rect 315500 664714 315528 685918
rect 316684 685908 316736 685914
rect 316684 685850 316736 685856
rect 295720 664686 296056 664714
rect 315376 664686 315528 664714
rect 305716 664006 306052 664034
rect 306024 662386 306052 664006
rect 316696 662386 316724 685850
rect 316788 665514 316816 686054
rect 345664 686044 345716 686050
rect 345664 685986 345716 685992
rect 361672 686044 361724 686050
rect 361672 685986 361724 685992
rect 371516 686044 371568 686050
rect 371516 685986 371568 685992
rect 389364 686044 389416 686050
rect 389364 685986 389416 685992
rect 399484 686044 399536 686050
rect 399484 685986 399536 685992
rect 333704 685976 333756 685982
rect 333704 685918 333756 685924
rect 333716 683876 333744 685918
rect 343364 685908 343416 685914
rect 343364 685850 343416 685856
rect 344284 685908 344336 685914
rect 344284 685850 344336 685856
rect 343376 683876 343404 685850
rect 323044 683318 324070 683346
rect 322846 674248 322902 674257
rect 322846 674183 322902 674192
rect 317418 673568 317474 673577
rect 317418 673503 317474 673512
rect 316776 665508 316828 665514
rect 316776 665450 316828 665456
rect 317432 665174 317460 673503
rect 322860 665174 322888 674183
rect 317420 665168 317472 665174
rect 317420 665110 317472 665116
rect 322848 665168 322900 665174
rect 322848 665110 322900 665116
rect 277676 662380 277728 662386
rect 277676 662322 277728 662328
rect 289084 662380 289136 662386
rect 289084 662322 289136 662328
rect 306012 662380 306064 662386
rect 306012 662322 306064 662328
rect 316684 662380 316736 662386
rect 316684 662322 316736 662328
rect 323044 662250 323072 683318
rect 323676 665508 323728 665514
rect 323676 665450 323728 665456
rect 323688 664714 323716 665450
rect 343548 665100 343600 665106
rect 343548 665042 343600 665048
rect 343560 664714 343588 665042
rect 323688 664686 324070 664714
rect 343390 664686 343588 664714
rect 333730 664006 333928 664034
rect 333900 662318 333928 664006
rect 344296 662318 344324 685850
rect 345020 683188 345072 683194
rect 345020 683130 345072 683136
rect 345032 673577 345060 683130
rect 345018 673568 345074 673577
rect 345018 673503 345074 673512
rect 345676 665106 345704 685986
rect 352012 685976 352064 685982
rect 352012 685918 352064 685924
rect 352024 683876 352052 685918
rect 361684 683876 361712 685986
rect 371332 685908 371384 685914
rect 371332 685850 371384 685856
rect 371344 683876 371372 685850
rect 350448 683188 350500 683194
rect 350448 683130 350500 683136
rect 350460 674257 350488 683130
rect 350446 674248 350502 674257
rect 350446 674183 350502 674192
rect 345664 665100 345716 665106
rect 345664 665042 345716 665048
rect 371528 664714 371556 685986
rect 374644 685976 374696 685982
rect 374644 685918 374696 685924
rect 373264 685908 373316 685914
rect 373264 685850 373316 685856
rect 371358 664686 371556 664714
rect 333888 662312 333940 662318
rect 333888 662254 333940 662260
rect 344284 662312 344336 662318
rect 344284 662254 344336 662260
rect 352024 662250 352052 664020
rect 361684 662386 361712 664020
rect 373276 662386 373304 685850
rect 373998 673568 374054 673577
rect 373998 673503 374054 673512
rect 374012 665174 374040 673503
rect 374000 665168 374052 665174
rect 374000 665110 374052 665116
rect 374656 662386 374684 685918
rect 389376 683890 389404 685986
rect 399024 685908 399076 685914
rect 399024 685850 399076 685856
rect 399036 683890 399064 685850
rect 389376 683862 389712 683890
rect 399036 683862 399372 683890
rect 379624 683318 380052 683346
rect 378048 683256 378100 683262
rect 378048 683198 378100 683204
rect 378060 674257 378088 683198
rect 378046 674248 378102 674257
rect 378046 674183 378102 674192
rect 361672 662380 361724 662386
rect 361672 662322 361724 662328
rect 373264 662380 373316 662386
rect 373264 662322 373316 662328
rect 374644 662380 374696 662386
rect 374644 662322 374696 662328
rect 379624 662318 379652 683318
rect 399496 664714 399524 685986
rect 400864 685908 400916 685914
rect 400864 685850 400916 685856
rect 399372 664686 399524 664714
rect 379716 664006 380052 664034
rect 389712 664006 390048 664034
rect 379716 662386 379744 664006
rect 379704 662380 379756 662386
rect 379704 662322 379756 662328
rect 390020 662318 390048 664006
rect 400876 662318 400904 685850
rect 408052 683876 408080 686054
rect 417700 686044 417752 686050
rect 417700 685986 417752 685992
rect 417712 683876 417740 685986
rect 428464 685976 428516 685982
rect 428464 685918 428516 685924
rect 427360 685908 427412 685914
rect 427360 685850 427412 685856
rect 427372 683876 427400 685850
rect 401600 683188 401652 683194
rect 401600 683130 401652 683136
rect 401612 673577 401640 683130
rect 405646 674248 405702 674257
rect 405646 674183 405702 674192
rect 401598 673568 401654 673577
rect 401598 673503 401654 673512
rect 405660 665174 405688 674183
rect 428476 673454 428504 685918
rect 428556 685908 428608 685914
rect 428556 685850 428608 685856
rect 427832 673426 428504 673454
rect 405648 665168 405700 665174
rect 405648 665110 405700 665116
rect 427832 664714 427860 673426
rect 427386 664686 427860 664714
rect 408052 662386 408080 664020
rect 408040 662380 408092 662386
rect 408040 662322 408092 662328
rect 417712 662318 417740 664020
rect 428568 662318 428596 685850
rect 428660 665854 428688 686054
rect 456156 686044 456208 686050
rect 456156 685986 456208 685992
rect 473360 686044 473412 686050
rect 473360 685986 473412 685992
rect 483480 686044 483532 686050
rect 483480 685986 483532 685992
rect 445668 685976 445720 685982
rect 445668 685918 445720 685924
rect 445680 683876 445708 685918
rect 455328 685908 455380 685914
rect 455328 685850 455380 685856
rect 456064 685908 456116 685914
rect 456064 685850 456116 685856
rect 455340 683876 455368 685850
rect 434824 683318 436034 683346
rect 429200 683256 429252 683262
rect 429200 683198 429252 683204
rect 429212 673577 429240 683198
rect 434628 683188 434680 683194
rect 434628 683130 434680 683136
rect 434640 674257 434668 683130
rect 434626 674248 434682 674257
rect 434626 674183 434682 674192
rect 429198 673568 429254 673577
rect 429198 673503 429254 673512
rect 428648 665848 428700 665854
rect 428648 665790 428700 665796
rect 379612 662312 379664 662318
rect 379612 662254 379664 662260
rect 390008 662312 390060 662318
rect 390008 662254 390060 662260
rect 400864 662312 400916 662318
rect 400864 662254 400916 662260
rect 417700 662312 417752 662318
rect 417700 662254 417752 662260
rect 428556 662312 428608 662318
rect 428556 662254 428608 662260
rect 434824 662250 434852 683318
rect 455696 668772 455748 668778
rect 455696 668714 455748 668720
rect 435732 665848 435784 665854
rect 435732 665790 435784 665796
rect 435744 664714 435772 665790
rect 455708 664714 455736 668714
rect 435744 664686 436034 664714
rect 455354 664686 455736 664714
rect 445680 662318 445708 664020
rect 456076 662318 456104 685850
rect 456168 668778 456196 685986
rect 464344 685976 464396 685982
rect 464344 685918 464396 685924
rect 464356 683890 464384 685918
rect 464048 683862 464384 683890
rect 473372 683890 473400 685986
rect 483020 685908 483072 685914
rect 483020 685850 483072 685856
rect 483032 683890 483060 685850
rect 473372 683862 473708 683890
rect 483032 683862 483368 683890
rect 462226 674248 462282 674257
rect 462226 674183 462282 674192
rect 458178 673568 458234 673577
rect 458178 673503 458234 673512
rect 456156 668772 456208 668778
rect 456156 668714 456208 668720
rect 458192 665174 458220 673503
rect 462240 665174 462268 674183
rect 458180 665168 458232 665174
rect 458180 665110 458232 665116
rect 462228 665168 462280 665174
rect 462228 665110 462280 665116
rect 483492 664714 483520 685986
rect 483664 685976 483716 685982
rect 483664 685918 483716 685924
rect 483676 665310 483704 685918
rect 485044 685908 485096 685914
rect 485044 685850 485096 685856
rect 483664 665304 483716 665310
rect 483664 665246 483716 665252
rect 483368 664686 483520 664714
rect 463804 664006 464048 664034
rect 473708 664006 474044 664034
rect 445668 662312 445720 662318
rect 445668 662254 445720 662260
rect 456064 662312 456116 662318
rect 456064 662254 456116 662260
rect 463804 662250 463832 664006
rect 474016 662386 474044 664006
rect 485056 662386 485084 685850
rect 485780 683188 485832 683194
rect 485780 683130 485832 683136
rect 489828 683188 489880 683194
rect 489828 683130 489880 683136
rect 485792 673577 485820 683130
rect 489840 674257 489868 683130
rect 489826 674248 489882 674257
rect 489826 674183 489882 674192
rect 485778 673568 485834 673577
rect 485778 673503 485834 673512
rect 474004 662380 474056 662386
rect 474004 662322 474056 662328
rect 485044 662380 485096 662386
rect 485044 662322 485096 662328
rect 238852 662244 238904 662250
rect 238852 662186 238904 662192
rect 268016 662244 268068 662250
rect 268016 662186 268068 662192
rect 323032 662244 323084 662250
rect 323032 662186 323084 662192
rect 352012 662244 352064 662250
rect 352012 662186 352064 662192
rect 434812 662244 434864 662250
rect 434812 662186 434864 662192
rect 463792 662244 463844 662250
rect 463792 662186 463844 662192
rect 296352 658504 296404 658510
rect 296352 658446 296404 658452
rect 316776 658504 316828 658510
rect 316776 658446 316828 658452
rect 408040 658504 408092 658510
rect 408040 658446 408092 658452
rect 428648 658504 428700 658510
rect 428648 658446 428700 658452
rect 260196 658436 260248 658442
rect 260196 658378 260248 658384
rect 277676 658436 277728 658442
rect 277676 658378 277728 658384
rect 287520 658436 287572 658442
rect 287520 658378 287572 658384
rect 249708 658368 249760 658374
rect 249708 658310 249760 658316
rect 249720 656948 249748 658310
rect 259368 658300 259420 658306
rect 259368 658242 259420 658248
rect 260104 658300 260156 658306
rect 260104 658242 260156 658248
rect 259380 656948 259408 658242
rect 238864 656254 240074 656282
rect 238668 655648 238720 655654
rect 238668 655590 238720 655596
rect 238680 647329 238708 655590
rect 238666 647320 238722 647329
rect 238666 647255 238722 647264
rect 238864 634642 238892 656254
rect 259736 640824 259788 640830
rect 259736 640766 259788 640772
rect 239772 639396 239824 639402
rect 239772 639338 239824 639344
rect 239784 637786 239812 639338
rect 259748 637786 259776 640766
rect 239784 637758 240074 637786
rect 259394 637758 259776 637786
rect 238852 634636 238904 634642
rect 238852 634578 238904 634584
rect 249720 634574 249748 637092
rect 260116 634574 260144 658242
rect 260208 640830 260236 658378
rect 268016 658368 268068 658374
rect 268016 658310 268068 658316
rect 268028 656948 268056 658310
rect 277688 656948 277716 658378
rect 287336 658300 287388 658306
rect 287336 658242 287388 658248
rect 287348 656948 287376 658242
rect 262220 655580 262272 655586
rect 262220 655522 262272 655528
rect 266268 655580 266320 655586
rect 266268 655522 266320 655528
rect 262232 646649 262260 655522
rect 266280 647329 266308 655522
rect 266266 647320 266322 647329
rect 266266 647255 266322 647264
rect 262218 646640 262274 646649
rect 262218 646575 262274 646584
rect 260196 640824 260248 640830
rect 260196 640766 260248 640772
rect 287532 637786 287560 658378
rect 287704 658368 287756 658374
rect 287704 658310 287756 658316
rect 287716 639810 287744 658310
rect 289084 658300 289136 658306
rect 289084 658242 289136 658248
rect 287704 639804 287756 639810
rect 287704 639746 287756 639752
rect 287362 637758 287560 637786
rect 268028 634642 268056 637092
rect 277688 634642 277716 637092
rect 289096 634642 289124 658242
rect 296364 656962 296392 658446
rect 305368 658436 305420 658442
rect 305368 658378 305420 658384
rect 296056 656934 296392 656962
rect 305380 656962 305408 658378
rect 315488 658368 315540 658374
rect 315488 658310 315540 658316
rect 315028 658300 315080 658306
rect 315028 658242 315080 658248
rect 315040 656962 315068 658242
rect 305380 656934 305716 656962
rect 315040 656934 315376 656962
rect 289820 655648 289872 655654
rect 289820 655590 289872 655596
rect 293868 655648 293920 655654
rect 293868 655590 293920 655596
rect 289832 646649 289860 655590
rect 293880 647329 293908 655590
rect 293866 647320 293922 647329
rect 293866 647255 293922 647264
rect 289818 646640 289874 646649
rect 289818 646575 289874 646584
rect 295708 639804 295760 639810
rect 295708 639746 295760 639752
rect 295720 637786 295748 639746
rect 315500 637786 315528 658310
rect 316684 658300 316736 658306
rect 316684 658242 316736 658248
rect 295720 637758 296056 637786
rect 315376 637758 315528 637786
rect 305716 637078 306052 637106
rect 306024 634642 306052 637078
rect 316696 634642 316724 658242
rect 316788 639402 316816 658446
rect 345664 658436 345716 658442
rect 345664 658378 345716 658384
rect 361672 658436 361724 658442
rect 361672 658378 361724 658384
rect 371516 658436 371568 658442
rect 371516 658378 371568 658384
rect 389364 658436 389416 658442
rect 389364 658378 389416 658384
rect 399484 658436 399536 658442
rect 399484 658378 399536 658384
rect 333704 658368 333756 658374
rect 333704 658310 333756 658316
rect 333716 656948 333744 658310
rect 343364 658300 343416 658306
rect 343364 658242 343416 658248
rect 344284 658300 344336 658306
rect 344284 658242 344336 658248
rect 343376 656948 343404 658242
rect 323044 656254 324070 656282
rect 317420 655580 317472 655586
rect 317420 655522 317472 655528
rect 322848 655580 322900 655586
rect 322848 655522 322900 655528
rect 317432 646649 317460 655522
rect 322860 647329 322888 655522
rect 322846 647320 322902 647329
rect 322846 647255 322902 647264
rect 317418 646640 317474 646649
rect 317418 646575 317474 646584
rect 316776 639396 316828 639402
rect 316776 639338 316828 639344
rect 323044 634642 323072 656254
rect 323676 639396 323728 639402
rect 323676 639338 323728 639344
rect 323688 637786 323716 639338
rect 323688 637758 324070 637786
rect 343640 637560 343692 637566
rect 343390 637508 343640 637514
rect 343390 637502 343692 637508
rect 343390 637486 343680 637502
rect 268016 634636 268068 634642
rect 268016 634578 268068 634584
rect 277676 634636 277728 634642
rect 277676 634578 277728 634584
rect 289084 634636 289136 634642
rect 289084 634578 289136 634584
rect 306012 634636 306064 634642
rect 306012 634578 306064 634584
rect 316684 634636 316736 634642
rect 316684 634578 316736 634584
rect 323032 634636 323084 634642
rect 323032 634578 323084 634584
rect 333716 634574 333744 637092
rect 344296 634574 344324 658242
rect 345020 655648 345072 655654
rect 345020 655590 345072 655596
rect 345032 646649 345060 655590
rect 345018 646640 345074 646649
rect 345018 646575 345074 646584
rect 345676 637566 345704 658378
rect 352012 658368 352064 658374
rect 352012 658310 352064 658316
rect 352024 656948 352052 658310
rect 361684 656948 361712 658378
rect 371332 658300 371384 658306
rect 371332 658242 371384 658248
rect 371344 656948 371372 658242
rect 350448 655648 350500 655654
rect 350448 655590 350500 655596
rect 350460 647329 350488 655590
rect 350446 647320 350502 647329
rect 350446 647255 350502 647264
rect 371528 637786 371556 658378
rect 374644 658368 374696 658374
rect 374644 658310 374696 658316
rect 373264 658300 373316 658306
rect 373264 658242 373316 658248
rect 371358 637758 371556 637786
rect 345664 637560 345716 637566
rect 345664 637502 345716 637508
rect 352024 634642 352052 637092
rect 361684 634642 361712 637092
rect 373276 634642 373304 658242
rect 374000 655580 374052 655586
rect 374000 655522 374052 655528
rect 374012 646649 374040 655522
rect 373998 646640 374054 646649
rect 373998 646575 374054 646584
rect 374656 634778 374684 658310
rect 389376 656962 389404 658378
rect 399024 658300 399076 658306
rect 399024 658242 399076 658248
rect 399036 656962 399064 658242
rect 389376 656934 389712 656962
rect 399036 656934 399372 656962
rect 379624 656254 380052 656282
rect 378048 655716 378100 655722
rect 378048 655658 378100 655664
rect 378060 647329 378088 655658
rect 378046 647320 378102 647329
rect 378046 647255 378102 647264
rect 374644 634772 374696 634778
rect 374644 634714 374696 634720
rect 379624 634642 379652 656254
rect 399496 637786 399524 658378
rect 400864 658300 400916 658306
rect 400864 658242 400916 658248
rect 399372 637758 399524 637786
rect 379716 637078 380052 637106
rect 389712 637078 390048 637106
rect 379716 634778 379744 637078
rect 379704 634772 379756 634778
rect 379704 634714 379756 634720
rect 352012 634636 352064 634642
rect 352012 634578 352064 634584
rect 361672 634636 361724 634642
rect 361672 634578 361724 634584
rect 373264 634636 373316 634642
rect 373264 634578 373316 634584
rect 379612 634636 379664 634642
rect 379612 634578 379664 634584
rect 390020 634574 390048 637078
rect 400876 634574 400904 658242
rect 408052 656948 408080 658446
rect 417700 658436 417752 658442
rect 417700 658378 417752 658384
rect 417712 656948 417740 658378
rect 428464 658368 428516 658374
rect 428464 658310 428516 658316
rect 427360 658300 427412 658306
rect 427360 658242 427412 658248
rect 427372 656948 427400 658242
rect 401600 655648 401652 655654
rect 401600 655590 401652 655596
rect 401612 646649 401640 655590
rect 405648 655580 405700 655586
rect 405648 655522 405700 655528
rect 405660 647329 405688 655522
rect 405646 647320 405702 647329
rect 405646 647255 405702 647264
rect 401598 646640 401654 646649
rect 401598 646575 401654 646584
rect 428476 644474 428504 658310
rect 428556 658300 428608 658306
rect 428556 658242 428608 658248
rect 427832 644446 428504 644474
rect 427832 637514 427860 644446
rect 427386 637486 427860 637514
rect 408052 634642 408080 637092
rect 417712 634642 417740 637092
rect 428568 634642 428596 658242
rect 428660 639606 428688 658446
rect 456064 658436 456116 658442
rect 456064 658378 456116 658384
rect 473360 658436 473412 658442
rect 473360 658378 473412 658384
rect 483480 658436 483532 658442
rect 483480 658378 483532 658384
rect 445668 658368 445720 658374
rect 445668 658310 445720 658316
rect 445680 656948 445708 658310
rect 455328 658300 455380 658306
rect 455328 658242 455380 658248
rect 455340 656948 455368 658242
rect 434824 656254 436034 656282
rect 429200 655716 429252 655722
rect 429200 655658 429252 655664
rect 429212 646649 429240 655658
rect 434628 655648 434680 655654
rect 434628 655590 434680 655596
rect 434640 647329 434668 655590
rect 434626 647320 434682 647329
rect 434626 647255 434682 647264
rect 429198 646640 429254 646649
rect 429198 646575 429254 646584
rect 428648 639600 428700 639606
rect 428648 639542 428700 639548
rect 434824 634642 434852 656254
rect 456076 644474 456104 658378
rect 464344 658368 464396 658374
rect 464344 658310 464396 658316
rect 456156 658300 456208 658306
rect 456156 658242 456208 658248
rect 455800 644446 456104 644474
rect 435732 639600 435784 639606
rect 435732 639542 435784 639548
rect 435744 637786 435772 639542
rect 455800 637786 455828 644446
rect 435744 637758 436034 637786
rect 455354 637758 455828 637786
rect 408040 634636 408092 634642
rect 408040 634578 408092 634584
rect 417700 634636 417752 634642
rect 417700 634578 417752 634584
rect 428556 634636 428608 634642
rect 428556 634578 428608 634584
rect 434812 634636 434864 634642
rect 434812 634578 434864 634584
rect 445680 634574 445708 637092
rect 456168 634574 456196 658242
rect 464356 656962 464384 658310
rect 464048 656934 464384 656962
rect 473372 656962 473400 658378
rect 483020 658300 483072 658306
rect 483020 658242 483072 658248
rect 483032 656962 483060 658242
rect 473372 656934 473708 656962
rect 483032 656934 483368 656962
rect 463700 655716 463752 655722
rect 463700 655658 463752 655664
rect 458180 655580 458232 655586
rect 458180 655522 458232 655528
rect 458192 646649 458220 655522
rect 463712 654090 463740 655658
rect 462228 654084 462280 654090
rect 462228 654026 462280 654032
rect 463700 654084 463752 654090
rect 463700 654026 463752 654032
rect 462240 647329 462268 654026
rect 462226 647320 462282 647329
rect 462226 647255 462282 647264
rect 458178 646640 458234 646649
rect 458178 646575 458234 646584
rect 483492 637786 483520 658378
rect 483664 658368 483716 658374
rect 483664 658310 483716 658316
rect 483676 639402 483704 658310
rect 485044 658300 485096 658306
rect 485044 658242 485096 658248
rect 483664 639396 483716 639402
rect 483664 639338 483716 639344
rect 483368 637758 483520 637786
rect 463804 637078 464048 637106
rect 473708 637078 474044 637106
rect 463804 634642 463832 637078
rect 474016 634642 474044 637078
rect 485056 634642 485084 658242
rect 485780 655648 485832 655654
rect 485780 655590 485832 655596
rect 485792 646649 485820 655590
rect 489828 655580 489880 655586
rect 489828 655522 489880 655528
rect 489840 647329 489868 655522
rect 489826 647320 489882 647329
rect 489826 647255 489882 647264
rect 485778 646640 485834 646649
rect 485778 646575 485834 646584
rect 463792 634636 463844 634642
rect 463792 634578 463844 634584
rect 474004 634636 474056 634642
rect 474004 634578 474056 634584
rect 485044 634636 485096 634642
rect 485044 634578 485096 634584
rect 249708 634568 249760 634574
rect 249708 634510 249760 634516
rect 260104 634568 260156 634574
rect 260104 634510 260156 634516
rect 333704 634568 333756 634574
rect 333704 634510 333756 634516
rect 344284 634568 344336 634574
rect 344284 634510 344336 634516
rect 390008 634568 390060 634574
rect 390008 634510 390060 634516
rect 400864 634568 400916 634574
rect 400864 634510 400916 634516
rect 445668 634568 445720 634574
rect 445668 634510 445720 634516
rect 456156 634568 456208 634574
rect 456156 634510 456208 634516
rect 408040 632324 408092 632330
rect 408040 632266 408092 632272
rect 428648 632324 428700 632330
rect 428648 632266 428700 632272
rect 260104 632256 260156 632262
rect 260104 632198 260156 632204
rect 277676 632256 277728 632262
rect 277676 632198 277728 632204
rect 287520 632256 287572 632262
rect 287520 632198 287572 632204
rect 305368 632256 305420 632262
rect 305368 632198 305420 632204
rect 315488 632256 315540 632262
rect 315488 632198 315540 632204
rect 333704 632256 333756 632262
rect 333704 632198 333756 632204
rect 345664 632256 345716 632262
rect 345664 632198 345716 632204
rect 361672 632256 361724 632262
rect 361672 632198 361724 632204
rect 371516 632256 371568 632262
rect 371516 632198 371568 632204
rect 389364 632256 389416 632262
rect 389364 632198 389416 632204
rect 399484 632256 399536 632262
rect 399484 632198 399536 632204
rect 249708 632188 249760 632194
rect 249708 632130 249760 632136
rect 249720 629884 249748 632130
rect 259368 632120 259420 632126
rect 259368 632062 259420 632068
rect 259380 629884 259408 632062
rect 238864 629326 240074 629354
rect 238666 620256 238722 620265
rect 238666 620191 238722 620200
rect 238680 611250 238708 620191
rect 238668 611244 238720 611250
rect 238668 611186 238720 611192
rect 238864 608462 238892 629326
rect 260116 615494 260144 632198
rect 268016 632188 268068 632194
rect 268016 632130 268068 632136
rect 260196 632120 260248 632126
rect 260196 632062 260248 632068
rect 259840 615466 260144 615494
rect 239772 611992 239824 611998
rect 239772 611934 239824 611940
rect 239784 610722 239812 611934
rect 259840 610722 259868 615466
rect 239784 610694 240074 610722
rect 259394 610694 259868 610722
rect 238852 608456 238904 608462
rect 238852 608398 238904 608404
rect 249720 608394 249748 610028
rect 260208 608394 260236 632062
rect 268028 629884 268056 632130
rect 277688 629884 277716 632198
rect 287336 632120 287388 632126
rect 287336 632062 287388 632068
rect 287348 629884 287376 632062
rect 266266 620256 266322 620265
rect 266266 620191 266322 620200
rect 262218 619576 262274 619585
rect 262218 619511 262274 619520
rect 262232 611318 262260 619511
rect 266280 611318 266308 620191
rect 262220 611312 262272 611318
rect 262220 611254 262272 611260
rect 266268 611312 266320 611318
rect 266268 611254 266320 611260
rect 287532 610722 287560 632198
rect 287704 632188 287756 632194
rect 287704 632130 287756 632136
rect 296352 632188 296404 632194
rect 296352 632130 296404 632136
rect 287716 611930 287744 632130
rect 289084 632120 289136 632126
rect 289084 632062 289136 632068
rect 287704 611924 287756 611930
rect 287704 611866 287756 611872
rect 287362 610694 287560 610722
rect 268028 608462 268056 610028
rect 277688 608462 277716 610028
rect 289096 608462 289124 632062
rect 296364 629898 296392 632130
rect 296056 629870 296392 629898
rect 305380 629898 305408 632198
rect 315028 632120 315080 632126
rect 315028 632062 315080 632068
rect 315040 629898 315068 632062
rect 305380 629870 305716 629898
rect 315040 629870 315376 629898
rect 293866 620256 293922 620265
rect 293866 620191 293922 620200
rect 289818 619576 289874 619585
rect 289818 619511 289874 619520
rect 289832 611250 289860 619511
rect 293880 611250 293908 620191
rect 295708 611924 295760 611930
rect 295708 611866 295760 611872
rect 289820 611244 289872 611250
rect 289820 611186 289872 611192
rect 293868 611244 293920 611250
rect 293868 611186 293920 611192
rect 295720 610722 295748 611866
rect 315500 610722 315528 632198
rect 316776 632188 316828 632194
rect 316776 632130 316828 632136
rect 316684 632120 316736 632126
rect 316684 632062 316736 632068
rect 295720 610694 296056 610722
rect 315376 610694 315528 610722
rect 305716 610014 306052 610042
rect 306024 608462 306052 610014
rect 316696 608462 316724 632062
rect 316788 612066 316816 632130
rect 333716 629884 333744 632198
rect 343364 632120 343416 632126
rect 343364 632062 343416 632068
rect 344284 632120 344336 632126
rect 344284 632062 344336 632068
rect 343376 629884 343404 632062
rect 323044 629326 324070 629354
rect 322846 620256 322902 620265
rect 322846 620191 322902 620200
rect 317418 619576 317474 619585
rect 317418 619511 317474 619520
rect 316776 612060 316828 612066
rect 316776 612002 316828 612008
rect 317432 611318 317460 619511
rect 322860 611318 322888 620191
rect 317420 611312 317472 611318
rect 317420 611254 317472 611260
rect 322848 611312 322900 611318
rect 322848 611254 322900 611260
rect 323044 608462 323072 629326
rect 323676 612060 323728 612066
rect 323676 612002 323728 612008
rect 323688 610722 323716 612002
rect 323688 610694 324070 610722
rect 268016 608456 268068 608462
rect 268016 608398 268068 608404
rect 277676 608456 277728 608462
rect 277676 608398 277728 608404
rect 289084 608456 289136 608462
rect 289084 608398 289136 608404
rect 306012 608456 306064 608462
rect 306012 608398 306064 608404
rect 316684 608456 316736 608462
rect 316684 608398 316736 608404
rect 323032 608456 323084 608462
rect 323032 608398 323084 608404
rect 333716 608394 333744 610028
rect 343376 608598 343404 610028
rect 343364 608592 343416 608598
rect 343364 608534 343416 608540
rect 344296 608394 344324 632062
rect 345018 619576 345074 619585
rect 345018 619511 345074 619520
rect 345032 611250 345060 619511
rect 345020 611244 345072 611250
rect 345020 611186 345072 611192
rect 345676 608598 345704 632198
rect 352012 632188 352064 632194
rect 352012 632130 352064 632136
rect 352024 629884 352052 632130
rect 361684 629884 361712 632198
rect 371332 632120 371384 632126
rect 371332 632062 371384 632068
rect 371344 629884 371372 632062
rect 350446 620256 350502 620265
rect 350446 620191 350502 620200
rect 350460 611250 350488 620191
rect 350448 611244 350500 611250
rect 350448 611186 350500 611192
rect 371528 610722 371556 632198
rect 374644 632188 374696 632194
rect 374644 632130 374696 632136
rect 373264 632120 373316 632126
rect 373264 632062 373316 632068
rect 371358 610694 371556 610722
rect 345664 608592 345716 608598
rect 345664 608534 345716 608540
rect 352024 608462 352052 610028
rect 361684 608462 361712 610028
rect 373276 608462 373304 632062
rect 373998 619576 374054 619585
rect 373998 619511 374054 619520
rect 374012 611318 374040 619511
rect 374000 611312 374052 611318
rect 374000 611254 374052 611260
rect 374656 608598 374684 632130
rect 389376 629898 389404 632198
rect 399024 632120 399076 632126
rect 399024 632062 399076 632068
rect 399036 629898 399064 632062
rect 389376 629870 389712 629898
rect 399036 629870 399372 629898
rect 379624 629326 380052 629354
rect 378046 620256 378102 620265
rect 378046 620191 378102 620200
rect 378060 611182 378088 620191
rect 378048 611176 378100 611182
rect 378048 611118 378100 611124
rect 374644 608592 374696 608598
rect 374644 608534 374696 608540
rect 379624 608462 379652 629326
rect 399496 610722 399524 632198
rect 400864 632120 400916 632126
rect 400864 632062 400916 632068
rect 399372 610694 399524 610722
rect 379716 610014 380052 610042
rect 389712 610014 390048 610042
rect 379716 608598 379744 610014
rect 379704 608592 379756 608598
rect 379704 608534 379756 608540
rect 352012 608456 352064 608462
rect 352012 608398 352064 608404
rect 361672 608456 361724 608462
rect 361672 608398 361724 608404
rect 373264 608456 373316 608462
rect 373264 608398 373316 608404
rect 379612 608456 379664 608462
rect 379612 608398 379664 608404
rect 390020 608394 390048 610014
rect 400876 608394 400904 632062
rect 408052 629884 408080 632266
rect 417700 632256 417752 632262
rect 417700 632198 417752 632204
rect 417712 629884 417740 632198
rect 428464 632188 428516 632194
rect 428464 632130 428516 632136
rect 427360 632120 427412 632126
rect 427360 632062 427412 632068
rect 427372 629884 427400 632062
rect 405646 620256 405702 620265
rect 405646 620191 405702 620200
rect 401598 619576 401654 619585
rect 401598 619511 401654 619520
rect 401612 611250 401640 619511
rect 405660 611318 405688 620191
rect 428476 615494 428504 632130
rect 428556 632120 428608 632126
rect 428556 632062 428608 632068
rect 427832 615466 428504 615494
rect 405648 611312 405700 611318
rect 405648 611254 405700 611260
rect 401600 611244 401652 611250
rect 401600 611186 401652 611192
rect 427832 610722 427860 615466
rect 427386 610694 427860 610722
rect 408052 608462 408080 610028
rect 417712 608462 417740 610028
rect 428568 608462 428596 632062
rect 428660 612066 428688 632266
rect 456156 632256 456208 632262
rect 456156 632198 456208 632204
rect 473360 632256 473412 632262
rect 473360 632198 473412 632204
rect 483480 632256 483532 632262
rect 483480 632198 483532 632204
rect 445668 632188 445720 632194
rect 445668 632130 445720 632136
rect 445680 629884 445708 632130
rect 455328 632120 455380 632126
rect 455328 632062 455380 632068
rect 456064 632120 456116 632126
rect 456064 632062 456116 632068
rect 455340 629884 455368 632062
rect 434824 629326 436034 629354
rect 434626 620256 434682 620265
rect 434626 620191 434682 620200
rect 429198 619576 429254 619585
rect 429198 619511 429254 619520
rect 428648 612060 428700 612066
rect 428648 612002 428700 612008
rect 429212 611182 429240 619511
rect 434640 611182 434668 620191
rect 429200 611176 429252 611182
rect 429200 611118 429252 611124
rect 434628 611176 434680 611182
rect 434628 611118 434680 611124
rect 434824 608462 434852 629326
rect 455696 612808 455748 612814
rect 455696 612750 455748 612756
rect 435732 612060 435784 612066
rect 435732 612002 435784 612008
rect 435744 610722 435772 612002
rect 455708 610722 455736 612750
rect 435744 610694 436034 610722
rect 455354 610694 455736 610722
rect 408040 608456 408092 608462
rect 408040 608398 408092 608404
rect 417700 608456 417752 608462
rect 417700 608398 417752 608404
rect 428556 608456 428608 608462
rect 428556 608398 428608 608404
rect 434812 608456 434864 608462
rect 434812 608398 434864 608404
rect 445680 608394 445708 610028
rect 456076 608394 456104 632062
rect 456168 612814 456196 632198
rect 464344 632188 464396 632194
rect 464344 632130 464396 632136
rect 464356 629898 464384 632130
rect 464048 629870 464384 629898
rect 473372 629898 473400 632198
rect 483020 632120 483072 632126
rect 483020 632062 483072 632068
rect 483032 629898 483060 632062
rect 473372 629870 473708 629898
rect 483032 629870 483368 629898
rect 462226 620256 462282 620265
rect 462226 620191 462282 620200
rect 458178 619576 458234 619585
rect 458178 619511 458234 619520
rect 456156 612808 456208 612814
rect 456156 612750 456208 612756
rect 458192 611318 458220 619511
rect 458180 611312 458232 611318
rect 458180 611254 458232 611260
rect 462240 611250 462268 620191
rect 462228 611244 462280 611250
rect 462228 611186 462280 611192
rect 483492 610722 483520 632198
rect 483664 632188 483716 632194
rect 483664 632130 483716 632136
rect 483676 611794 483704 632130
rect 485044 632120 485096 632126
rect 485044 632062 485096 632068
rect 483664 611788 483716 611794
rect 483664 611730 483716 611736
rect 483368 610694 483520 610722
rect 463712 610014 464048 610042
rect 473708 610014 474044 610042
rect 463712 608462 463740 610014
rect 474016 608462 474044 610014
rect 485056 608462 485084 632062
rect 489826 620256 489882 620265
rect 489826 620191 489882 620200
rect 485778 619576 485834 619585
rect 485778 619511 485834 619520
rect 485792 611182 485820 619511
rect 489840 611318 489868 620191
rect 489828 611312 489880 611318
rect 489828 611254 489880 611260
rect 485780 611176 485832 611182
rect 485780 611118 485832 611124
rect 463700 608456 463752 608462
rect 463700 608398 463752 608404
rect 474004 608456 474056 608462
rect 474004 608398 474056 608404
rect 485044 608456 485096 608462
rect 485044 608398 485096 608404
rect 249708 608388 249760 608394
rect 249708 608330 249760 608336
rect 260196 608388 260248 608394
rect 260196 608330 260248 608336
rect 333704 608388 333756 608394
rect 333704 608330 333756 608336
rect 344284 608388 344336 608394
rect 344284 608330 344336 608336
rect 390008 608388 390060 608394
rect 390008 608330 390060 608336
rect 400864 608388 400916 608394
rect 400864 608330 400916 608336
rect 445668 608388 445720 608394
rect 445668 608330 445720 608336
rect 456064 608388 456116 608394
rect 456064 608330 456116 608336
rect 261484 604784 261536 604790
rect 261484 604726 261536 604732
rect 249708 604648 249760 604654
rect 249708 604590 249760 604596
rect 260196 604648 260248 604654
rect 260196 604590 260248 604596
rect 249720 602956 249748 604590
rect 259368 604580 259420 604586
rect 259368 604522 259420 604528
rect 259380 602956 259408 604522
rect 260104 604512 260156 604518
rect 260104 604454 260156 604460
rect 238864 602262 240074 602290
rect 238666 593328 238722 593337
rect 238666 593263 238722 593272
rect 238680 583642 238708 593263
rect 238668 583636 238720 583642
rect 238668 583578 238720 583584
rect 238864 580854 238892 602262
rect 259736 584792 259788 584798
rect 259736 584734 259788 584740
rect 239772 584452 239824 584458
rect 239772 584394 239824 584400
rect 239784 583794 239812 584394
rect 259748 583794 259776 584734
rect 239784 583766 240074 583794
rect 259394 583766 259776 583794
rect 238852 580848 238904 580854
rect 238852 580790 238904 580796
rect 249720 580786 249748 583100
rect 260116 580786 260144 604454
rect 260208 584798 260236 604590
rect 260196 584792 260248 584798
rect 260196 584734 260248 584740
rect 249708 580780 249760 580786
rect 249708 580722 249760 580728
rect 260104 580780 260156 580786
rect 260104 580722 260156 580728
rect 249708 578400 249760 578406
rect 249708 578342 249760 578348
rect 260196 578400 260248 578406
rect 260196 578342 260248 578348
rect 249720 575892 249748 578342
rect 259368 578264 259420 578270
rect 259368 578206 259420 578212
rect 260104 578264 260156 578270
rect 260104 578206 260156 578212
rect 259380 575892 259408 578206
rect 238864 575334 240074 575362
rect 238666 566264 238722 566273
rect 238666 566199 238722 566208
rect 238680 557462 238708 566199
rect 238668 557456 238720 557462
rect 238668 557398 238720 557404
rect 238864 554606 238892 575334
rect 259736 562352 259788 562358
rect 259736 562294 259788 562300
rect 239772 558204 239824 558210
rect 239772 558146 239824 558152
rect 239784 556730 239812 558146
rect 259748 556730 259776 562294
rect 239784 556702 240074 556730
rect 259394 556702 259776 556730
rect 249720 554674 249748 556036
rect 260116 554674 260144 578206
rect 260208 562358 260236 578342
rect 260196 562352 260248 562358
rect 260196 562294 260248 562300
rect 261496 554674 261524 604726
rect 408040 604716 408092 604722
rect 408040 604658 408092 604664
rect 428648 604716 428700 604722
rect 428648 604658 428700 604664
rect 277676 604648 277728 604654
rect 277676 604590 277728 604596
rect 287520 604648 287572 604654
rect 287520 604590 287572 604596
rect 305368 604648 305420 604654
rect 305368 604590 305420 604596
rect 315488 604648 315540 604654
rect 315488 604590 315540 604596
rect 333704 604648 333756 604654
rect 333704 604590 333756 604596
rect 345664 604648 345716 604654
rect 345664 604590 345716 604596
rect 361672 604648 361724 604654
rect 361672 604590 361724 604596
rect 371516 604648 371568 604654
rect 371516 604590 371568 604596
rect 389364 604648 389416 604654
rect 389364 604590 389416 604596
rect 399484 604648 399536 604654
rect 399484 604590 399536 604596
rect 268016 604580 268068 604586
rect 268016 604522 268068 604528
rect 268028 602956 268056 604522
rect 277688 602956 277716 604590
rect 287336 604512 287388 604518
rect 287336 604454 287388 604460
rect 287348 602956 287376 604454
rect 266266 593328 266322 593337
rect 266266 593263 266322 593272
rect 262218 592648 262274 592657
rect 262218 592583 262274 592592
rect 262232 583710 262260 592583
rect 266280 583710 266308 593263
rect 287532 583794 287560 604590
rect 287704 604580 287756 604586
rect 287704 604522 287756 604528
rect 296352 604580 296404 604586
rect 296352 604522 296404 604528
rect 287716 584186 287744 604522
rect 289084 604512 289136 604518
rect 289084 604454 289136 604460
rect 287704 584180 287756 584186
rect 287704 584122 287756 584128
rect 287362 583766 287560 583794
rect 262220 583704 262272 583710
rect 262220 583646 262272 583652
rect 266268 583704 266320 583710
rect 266268 583646 266320 583652
rect 268028 580854 268056 583100
rect 277688 580854 277716 583100
rect 289096 580854 289124 604454
rect 296364 602970 296392 604522
rect 296056 602942 296392 602970
rect 305380 602970 305408 604590
rect 315028 604512 315080 604518
rect 315028 604454 315080 604460
rect 315040 602970 315068 604454
rect 305380 602942 305716 602970
rect 315040 602942 315376 602970
rect 293866 593328 293922 593337
rect 293866 593263 293922 593272
rect 289818 592648 289874 592657
rect 289818 592583 289874 592592
rect 289832 583642 289860 592583
rect 293880 583642 293908 593263
rect 295708 584180 295760 584186
rect 295708 584122 295760 584128
rect 295720 583794 295748 584122
rect 315500 583794 315528 604590
rect 316776 604580 316828 604586
rect 316776 604522 316828 604528
rect 316684 604512 316736 604518
rect 316684 604454 316736 604460
rect 295720 583766 296056 583794
rect 315376 583766 315528 583794
rect 289820 583636 289872 583642
rect 289820 583578 289872 583584
rect 293868 583636 293920 583642
rect 293868 583578 293920 583584
rect 305716 583086 306052 583114
rect 306024 580854 306052 583086
rect 316696 580854 316724 604454
rect 316788 584322 316816 604522
rect 333716 602956 333744 604590
rect 343364 604512 343416 604518
rect 343364 604454 343416 604460
rect 344284 604512 344336 604518
rect 344284 604454 344336 604460
rect 343376 602956 343404 604454
rect 323044 602262 324070 602290
rect 322846 593328 322902 593337
rect 322846 593263 322902 593272
rect 317418 592648 317474 592657
rect 317418 592583 317474 592592
rect 316776 584316 316828 584322
rect 316776 584258 316828 584264
rect 317432 583710 317460 592583
rect 322860 583710 322888 593263
rect 317420 583704 317472 583710
rect 317420 583646 317472 583652
rect 322848 583704 322900 583710
rect 322848 583646 322900 583652
rect 323044 580854 323072 602262
rect 323860 584316 323912 584322
rect 323860 584258 323912 584264
rect 323872 583794 323900 584258
rect 323872 583766 324070 583794
rect 343390 583642 343680 583658
rect 343390 583636 343692 583642
rect 343390 583630 343640 583636
rect 343640 583578 343692 583584
rect 268016 580848 268068 580854
rect 268016 580790 268068 580796
rect 277676 580848 277728 580854
rect 277676 580790 277728 580796
rect 289084 580848 289136 580854
rect 289084 580790 289136 580796
rect 306012 580848 306064 580854
rect 306012 580790 306064 580796
rect 316684 580848 316736 580854
rect 316684 580790 316736 580796
rect 323032 580848 323084 580854
rect 323032 580790 323084 580796
rect 333716 580786 333744 583100
rect 344296 580786 344324 604454
rect 345018 592648 345074 592657
rect 345018 592583 345074 592592
rect 345032 583574 345060 592583
rect 345676 583642 345704 604590
rect 352012 604580 352064 604586
rect 352012 604522 352064 604528
rect 352024 602956 352052 604522
rect 361684 602956 361712 604590
rect 371332 604512 371384 604518
rect 371332 604454 371384 604460
rect 371344 602956 371372 604454
rect 350446 593328 350502 593337
rect 350446 593263 350502 593272
rect 350460 583642 350488 593263
rect 371528 583794 371556 604590
rect 374644 604580 374696 604586
rect 374644 604522 374696 604528
rect 373264 604512 373316 604518
rect 373264 604454 373316 604460
rect 371358 583766 371556 583794
rect 345664 583636 345716 583642
rect 345664 583578 345716 583584
rect 350448 583636 350500 583642
rect 350448 583578 350500 583584
rect 345020 583568 345072 583574
rect 345020 583510 345072 583516
rect 352024 580854 352052 583100
rect 361684 580854 361712 583100
rect 373276 580854 373304 604454
rect 373998 592648 374054 592657
rect 373998 592583 374054 592592
rect 374012 583710 374040 592583
rect 374000 583704 374052 583710
rect 374000 583646 374052 583652
rect 374656 580990 374684 604522
rect 389376 602970 389404 604590
rect 399024 604512 399076 604518
rect 399024 604454 399076 604460
rect 399036 602970 399064 604454
rect 389376 602942 389712 602970
rect 399036 602942 399372 602970
rect 379624 602262 380052 602290
rect 378046 593328 378102 593337
rect 378046 593263 378102 593272
rect 378060 583574 378088 593263
rect 378048 583568 378100 583574
rect 378048 583510 378100 583516
rect 374644 580984 374696 580990
rect 374644 580926 374696 580932
rect 379624 580854 379652 602262
rect 399496 583794 399524 604590
rect 400864 604512 400916 604518
rect 400864 604454 400916 604460
rect 399372 583766 399524 583794
rect 379716 583086 380052 583114
rect 389712 583086 390048 583114
rect 379716 580990 379744 583086
rect 379704 580984 379756 580990
rect 379704 580926 379756 580932
rect 352012 580848 352064 580854
rect 352012 580790 352064 580796
rect 361672 580848 361724 580854
rect 361672 580790 361724 580796
rect 373264 580848 373316 580854
rect 373264 580790 373316 580796
rect 379612 580848 379664 580854
rect 379612 580790 379664 580796
rect 390020 580786 390048 583086
rect 400876 580786 400904 604454
rect 408052 602956 408080 604658
rect 417700 604648 417752 604654
rect 417700 604590 417752 604596
rect 417712 602956 417740 604590
rect 428556 604580 428608 604586
rect 428556 604522 428608 604528
rect 427360 604512 427412 604518
rect 427360 604454 427412 604460
rect 428464 604512 428516 604518
rect 428464 604454 428516 604460
rect 427372 602956 427400 604454
rect 405646 593328 405702 593337
rect 405646 593263 405702 593272
rect 401598 592648 401654 592657
rect 401598 592583 401654 592592
rect 401612 583642 401640 592583
rect 405660 583710 405688 593263
rect 405648 583704 405700 583710
rect 405648 583646 405700 583652
rect 427386 583642 427768 583658
rect 401600 583636 401652 583642
rect 427386 583636 427780 583642
rect 427386 583630 427728 583636
rect 401600 583578 401652 583584
rect 427728 583578 427780 583584
rect 408052 580854 408080 583100
rect 417712 580854 417740 583100
rect 428476 580854 428504 604454
rect 428568 583642 428596 604522
rect 428660 584458 428688 604658
rect 456064 604648 456116 604654
rect 456064 604590 456116 604596
rect 473360 604648 473412 604654
rect 473360 604590 473412 604596
rect 483480 604648 483532 604654
rect 483480 604590 483532 604596
rect 445668 604580 445720 604586
rect 445668 604522 445720 604528
rect 445680 602956 445708 604522
rect 455328 604512 455380 604518
rect 455328 604454 455380 604460
rect 455340 602956 455368 604454
rect 434824 602262 436034 602290
rect 434626 593328 434682 593337
rect 434626 593263 434682 593272
rect 429198 592648 429254 592657
rect 429198 592583 429254 592592
rect 428648 584452 428700 584458
rect 428648 584394 428700 584400
rect 428556 583636 428608 583642
rect 428556 583578 428608 583584
rect 429212 583574 429240 592583
rect 434640 583642 434668 593263
rect 434628 583636 434680 583642
rect 434628 583578 434680 583584
rect 429200 583568 429252 583574
rect 429200 583510 429252 583516
rect 434824 580854 434852 602262
rect 456076 586514 456104 604590
rect 464344 604580 464396 604586
rect 464344 604522 464396 604528
rect 456156 604512 456208 604518
rect 456156 604454 456208 604460
rect 455800 586486 456104 586514
rect 435732 584452 435784 584458
rect 435732 584394 435784 584400
rect 435744 583794 435772 584394
rect 455800 583794 455828 586486
rect 435744 583766 436034 583794
rect 455354 583766 455828 583794
rect 408040 580848 408092 580854
rect 408040 580790 408092 580796
rect 417700 580848 417752 580854
rect 417700 580790 417752 580796
rect 428464 580848 428516 580854
rect 428464 580790 428516 580796
rect 434812 580848 434864 580854
rect 434812 580790 434864 580796
rect 445680 580786 445708 583100
rect 456168 580786 456196 604454
rect 464356 602970 464384 604522
rect 464048 602942 464384 602970
rect 473372 602970 473400 604590
rect 483020 604512 483072 604518
rect 483020 604454 483072 604460
rect 483032 602970 483060 604454
rect 473372 602942 473708 602970
rect 483032 602942 483368 602970
rect 462226 593328 462282 593337
rect 462226 593263 462282 593272
rect 458178 592648 458234 592657
rect 458178 592583 458234 592592
rect 458192 583710 458220 592583
rect 458180 583704 458232 583710
rect 458180 583646 458232 583652
rect 462240 583574 462268 593263
rect 483492 583794 483520 604590
rect 483664 604580 483716 604586
rect 483664 604522 483716 604528
rect 483676 584186 483704 604522
rect 485044 604512 485096 604518
rect 485044 604454 485096 604460
rect 483664 584180 483716 584186
rect 483664 584122 483716 584128
rect 483368 583766 483520 583794
rect 462228 583568 462280 583574
rect 462228 583510 462280 583516
rect 463712 583086 464048 583114
rect 473708 583086 474044 583114
rect 463712 580854 463740 583086
rect 474016 580854 474044 583086
rect 485056 580854 485084 604454
rect 489826 593328 489882 593337
rect 489826 593263 489882 593272
rect 485778 592648 485834 592657
rect 485778 592583 485834 592592
rect 485792 583642 485820 592583
rect 489840 583710 489868 593263
rect 489828 583704 489880 583710
rect 489828 583646 489880 583652
rect 485780 583636 485832 583642
rect 485780 583578 485832 583584
rect 463700 580848 463752 580854
rect 463700 580790 463752 580796
rect 474004 580848 474056 580854
rect 474004 580790 474056 580796
rect 485044 580848 485096 580854
rect 485044 580790 485096 580796
rect 333704 580780 333756 580786
rect 333704 580722 333756 580728
rect 344284 580780 344336 580786
rect 344284 580722 344336 580728
rect 390008 580780 390060 580786
rect 390008 580722 390060 580728
rect 400864 580780 400916 580786
rect 400864 580722 400916 580728
rect 445668 580780 445720 580786
rect 445668 580722 445720 580728
rect 456156 580780 456208 580786
rect 456156 580722 456208 580728
rect 296352 578468 296404 578474
rect 296352 578410 296404 578416
rect 316776 578468 316828 578474
rect 316776 578410 316828 578416
rect 408040 578468 408092 578474
rect 408040 578410 408092 578416
rect 428648 578468 428700 578474
rect 428648 578410 428700 578416
rect 277676 578400 277728 578406
rect 277676 578342 277728 578348
rect 287520 578400 287572 578406
rect 287520 578342 287572 578348
rect 268016 578332 268068 578338
rect 268016 578274 268068 578280
rect 268028 575892 268056 578274
rect 277688 575892 277716 578342
rect 287336 578264 287388 578270
rect 287336 578206 287388 578212
rect 287348 575892 287376 578206
rect 266266 566264 266322 566273
rect 266266 566199 266322 566208
rect 262218 565584 262274 565593
rect 262218 565519 262274 565528
rect 262232 557530 262260 565519
rect 266280 557530 266308 566199
rect 262220 557524 262272 557530
rect 262220 557466 262272 557472
rect 266268 557524 266320 557530
rect 266268 557466 266320 557472
rect 287532 556730 287560 578342
rect 287704 578332 287756 578338
rect 287704 578274 287756 578280
rect 287716 558890 287744 578274
rect 289084 578264 289136 578270
rect 289084 578206 289136 578212
rect 287704 558884 287756 558890
rect 287704 558826 287756 558832
rect 287362 556702 287560 556730
rect 249708 554668 249760 554674
rect 249708 554610 249760 554616
rect 260104 554668 260156 554674
rect 260104 554610 260156 554616
rect 261484 554668 261536 554674
rect 261484 554610 261536 554616
rect 268028 554606 268056 556036
rect 277688 554606 277716 556036
rect 289096 554606 289124 578206
rect 296364 575906 296392 578410
rect 305368 578400 305420 578406
rect 305368 578342 305420 578348
rect 296056 575878 296392 575906
rect 305380 575906 305408 578342
rect 315488 578332 315540 578338
rect 315488 578274 315540 578280
rect 315028 578264 315080 578270
rect 315028 578206 315080 578212
rect 315040 575906 315068 578206
rect 305380 575878 305716 575906
rect 315040 575878 315376 575906
rect 293866 566264 293922 566273
rect 293866 566199 293922 566208
rect 289818 565584 289874 565593
rect 289818 565519 289874 565528
rect 289832 557462 289860 565519
rect 293880 557462 293908 566199
rect 295708 558884 295760 558890
rect 295708 558826 295760 558832
rect 289820 557456 289872 557462
rect 289820 557398 289872 557404
rect 293868 557456 293920 557462
rect 293868 557398 293920 557404
rect 295720 556730 295748 558826
rect 315500 556730 315528 578274
rect 316684 578264 316736 578270
rect 316684 578206 316736 578212
rect 295720 556702 296056 556730
rect 315376 556702 315528 556730
rect 305716 556022 306052 556050
rect 306024 554606 306052 556022
rect 316696 554606 316724 578206
rect 316788 558890 316816 578410
rect 345664 578400 345716 578406
rect 345664 578342 345716 578348
rect 361672 578400 361724 578406
rect 361672 578342 361724 578348
rect 371516 578400 371568 578406
rect 371516 578342 371568 578348
rect 389364 578400 389416 578406
rect 389364 578342 389416 578348
rect 399484 578400 399536 578406
rect 399484 578342 399536 578348
rect 333704 578332 333756 578338
rect 333704 578274 333756 578280
rect 333716 575892 333744 578274
rect 343364 578264 343416 578270
rect 343364 578206 343416 578212
rect 344284 578264 344336 578270
rect 344284 578206 344336 578212
rect 343376 575892 343404 578206
rect 323044 575334 324070 575362
rect 322846 566264 322902 566273
rect 322846 566199 322902 566208
rect 317418 565584 317474 565593
rect 317418 565519 317474 565528
rect 316776 558884 316828 558890
rect 316776 558826 316828 558832
rect 317432 557530 317460 565519
rect 322860 557530 322888 566199
rect 317420 557524 317472 557530
rect 317420 557466 317472 557472
rect 322848 557524 322900 557530
rect 322848 557466 322900 557472
rect 323044 554606 323072 575334
rect 323676 558884 323728 558890
rect 323676 558826 323728 558832
rect 323688 556730 323716 558826
rect 343548 557456 343600 557462
rect 343548 557398 343600 557404
rect 343560 556730 343588 557398
rect 323688 556702 324070 556730
rect 343390 556702 343588 556730
rect 238852 554600 238904 554606
rect 238852 554542 238904 554548
rect 268016 554600 268068 554606
rect 268016 554542 268068 554548
rect 277676 554600 277728 554606
rect 277676 554542 277728 554548
rect 289084 554600 289136 554606
rect 289084 554542 289136 554548
rect 306012 554600 306064 554606
rect 306012 554542 306064 554548
rect 316684 554600 316736 554606
rect 316684 554542 316736 554548
rect 323032 554600 323084 554606
rect 323032 554542 323084 554548
rect 333716 554538 333744 556036
rect 344296 554538 344324 578206
rect 345018 565584 345074 565593
rect 345018 565519 345074 565528
rect 345032 557394 345060 565519
rect 345676 557462 345704 578342
rect 352012 578332 352064 578338
rect 352012 578274 352064 578280
rect 352024 575892 352052 578274
rect 361684 575892 361712 578342
rect 371332 578264 371384 578270
rect 371332 578206 371384 578212
rect 371344 575892 371372 578206
rect 350446 566264 350502 566273
rect 350446 566199 350502 566208
rect 350460 557462 350488 566199
rect 345664 557456 345716 557462
rect 345664 557398 345716 557404
rect 350448 557456 350500 557462
rect 350448 557398 350500 557404
rect 345020 557388 345072 557394
rect 345020 557330 345072 557336
rect 371528 556730 371556 578342
rect 374644 578332 374696 578338
rect 374644 578274 374696 578280
rect 373264 578264 373316 578270
rect 373264 578206 373316 578212
rect 371358 556702 371556 556730
rect 352024 554606 352052 556036
rect 361684 554606 361712 556036
rect 373276 554606 373304 578206
rect 373998 565584 374054 565593
rect 373998 565519 374054 565528
rect 374012 557530 374040 565519
rect 374000 557524 374052 557530
rect 374000 557466 374052 557472
rect 374656 554742 374684 578274
rect 389376 575906 389404 578342
rect 399024 578264 399076 578270
rect 399024 578206 399076 578212
rect 399036 575906 399064 578206
rect 389376 575878 389712 575906
rect 399036 575878 399372 575906
rect 379624 575334 380052 575362
rect 378046 566264 378102 566273
rect 378046 566199 378102 566208
rect 378060 557394 378088 566199
rect 378048 557388 378100 557394
rect 378048 557330 378100 557336
rect 374644 554736 374696 554742
rect 374644 554678 374696 554684
rect 379624 554606 379652 575334
rect 399496 556730 399524 578342
rect 400864 578264 400916 578270
rect 400864 578206 400916 578212
rect 399372 556702 399524 556730
rect 379716 556022 380052 556050
rect 389712 556022 390048 556050
rect 379716 554742 379744 556022
rect 379704 554736 379756 554742
rect 379704 554678 379756 554684
rect 352012 554600 352064 554606
rect 352012 554542 352064 554548
rect 361672 554600 361724 554606
rect 361672 554542 361724 554548
rect 373264 554600 373316 554606
rect 373264 554542 373316 554548
rect 379612 554600 379664 554606
rect 379612 554542 379664 554548
rect 390020 554538 390048 556022
rect 400876 554538 400904 578206
rect 408052 575892 408080 578410
rect 417700 578400 417752 578406
rect 417700 578342 417752 578348
rect 417712 575892 417740 578342
rect 428464 578332 428516 578338
rect 428464 578274 428516 578280
rect 427360 578264 427412 578270
rect 427360 578206 427412 578212
rect 427372 575892 427400 578206
rect 405646 566264 405702 566273
rect 405646 566199 405702 566208
rect 401598 565584 401654 565593
rect 401598 565519 401654 565528
rect 401612 557462 401640 565519
rect 405660 557530 405688 566199
rect 428476 557534 428504 578274
rect 428556 578264 428608 578270
rect 428556 578206 428608 578212
rect 405648 557524 405700 557530
rect 405648 557466 405700 557472
rect 427832 557506 428504 557534
rect 401600 557456 401652 557462
rect 401600 557398 401652 557404
rect 427832 556730 427860 557506
rect 427386 556702 427860 556730
rect 408052 554606 408080 556036
rect 417712 554606 417740 556036
rect 428568 554606 428596 578206
rect 428660 558210 428688 578410
rect 456156 578400 456208 578406
rect 456156 578342 456208 578348
rect 473544 578400 473596 578406
rect 473544 578342 473596 578348
rect 483480 578400 483532 578406
rect 483480 578342 483532 578348
rect 445668 578332 445720 578338
rect 445668 578274 445720 578280
rect 445680 575892 445708 578274
rect 455328 578264 455380 578270
rect 455328 578206 455380 578212
rect 456064 578264 456116 578270
rect 456064 578206 456116 578212
rect 455340 575892 455368 578206
rect 434824 575334 436034 575362
rect 434626 566264 434682 566273
rect 434626 566199 434682 566208
rect 429198 565584 429254 565593
rect 429198 565519 429254 565528
rect 428648 558204 428700 558210
rect 428648 558146 428700 558152
rect 429212 557394 429240 565519
rect 434640 557462 434668 566199
rect 434628 557456 434680 557462
rect 434628 557398 434680 557404
rect 429200 557388 429252 557394
rect 429200 557330 429252 557336
rect 434824 554606 434852 575334
rect 455696 562352 455748 562358
rect 455696 562294 455748 562300
rect 435732 558204 435784 558210
rect 435732 558146 435784 558152
rect 435744 556730 435772 558146
rect 455708 556730 455736 562294
rect 435744 556702 436034 556730
rect 455354 556702 455736 556730
rect 408040 554600 408092 554606
rect 408040 554542 408092 554548
rect 417700 554600 417752 554606
rect 417700 554542 417752 554548
rect 428556 554600 428608 554606
rect 428556 554542 428608 554548
rect 434812 554600 434864 554606
rect 434812 554542 434864 554548
rect 445680 554538 445708 556036
rect 456076 554538 456104 578206
rect 456168 562358 456196 578342
rect 464344 578332 464396 578338
rect 464344 578274 464396 578280
rect 464356 575906 464384 578274
rect 464048 575878 464384 575906
rect 473556 575906 473584 578342
rect 483204 578264 483256 578270
rect 483204 578206 483256 578212
rect 483216 575906 483244 578206
rect 473556 575878 473708 575906
rect 483216 575878 483368 575906
rect 462226 566264 462282 566273
rect 462226 566199 462282 566208
rect 458178 565584 458234 565593
rect 458178 565519 458234 565528
rect 456156 562352 456208 562358
rect 456156 562294 456208 562300
rect 458192 557530 458220 565519
rect 458180 557524 458232 557530
rect 458180 557466 458232 557472
rect 462240 557394 462268 566199
rect 462228 557388 462280 557394
rect 462228 557330 462280 557336
rect 483492 556730 483520 578342
rect 483664 578332 483716 578338
rect 483664 578274 483716 578280
rect 483676 558210 483704 578274
rect 485044 578264 485096 578270
rect 485044 578206 485096 578212
rect 483664 558204 483716 558210
rect 483664 558146 483716 558152
rect 483368 556702 483520 556730
rect 463712 556022 464048 556050
rect 473708 556022 474044 556050
rect 463712 554606 463740 556022
rect 474016 554606 474044 556022
rect 485056 554606 485084 578206
rect 489826 566264 489882 566273
rect 489826 566199 489882 566208
rect 485778 565584 485834 565593
rect 485778 565519 485834 565528
rect 485792 557462 485820 565519
rect 489840 557530 489868 566199
rect 489828 557524 489880 557530
rect 489828 557466 489880 557472
rect 485780 557456 485832 557462
rect 485780 557398 485832 557404
rect 463700 554600 463752 554606
rect 463700 554542 463752 554548
rect 474004 554600 474056 554606
rect 474004 554542 474056 554548
rect 485044 554600 485096 554606
rect 485044 554542 485096 554548
rect 333704 554532 333756 554538
rect 333704 554474 333756 554480
rect 344284 554532 344336 554538
rect 344284 554474 344336 554480
rect 390008 554532 390060 554538
rect 390008 554474 390060 554480
rect 400864 554532 400916 554538
rect 400864 554474 400916 554480
rect 445668 554532 445720 554538
rect 445668 554474 445720 554480
rect 456064 554532 456116 554538
rect 456064 554474 456116 554480
rect 261484 550928 261536 550934
rect 261484 550870 261536 550876
rect 249708 550792 249760 550798
rect 249708 550734 249760 550740
rect 260104 550792 260156 550798
rect 260104 550734 260156 550740
rect 249720 548964 249748 550734
rect 259368 550724 259420 550730
rect 259368 550666 259420 550672
rect 259380 548964 259408 550666
rect 238864 548270 240074 548298
rect 238666 539336 238722 539345
rect 238666 539271 238722 539280
rect 238680 529854 238708 539271
rect 238668 529848 238720 529854
rect 238668 529790 238720 529796
rect 238864 526998 238892 548270
rect 260116 538214 260144 550734
rect 260196 550656 260248 550662
rect 260196 550598 260248 550604
rect 259840 538186 260144 538214
rect 239772 530256 239824 530262
rect 239772 530198 239824 530204
rect 239784 529666 239812 530198
rect 259840 529666 259868 538186
rect 239784 529638 240074 529666
rect 259394 529638 259868 529666
rect 238852 526992 238904 526998
rect 238852 526934 238904 526940
rect 249720 526930 249748 529108
rect 260208 526930 260236 550598
rect 249708 526924 249760 526930
rect 249708 526866 249760 526872
rect 260196 526924 260248 526930
rect 260196 526866 260248 526872
rect 260196 523184 260248 523190
rect 260196 523126 260248 523132
rect 249708 523116 249760 523122
rect 249708 523058 249760 523064
rect 249720 521900 249748 523058
rect 259368 523048 259420 523054
rect 259368 522990 259420 522996
rect 260104 523048 260156 523054
rect 260104 522990 260156 522996
rect 259380 521900 259408 522990
rect 238864 521206 240074 521234
rect 238668 520396 238720 520402
rect 238668 520338 238720 520344
rect 238680 512281 238708 520338
rect 238666 512272 238722 512281
rect 238666 512207 238722 512216
rect 238864 500818 238892 521206
rect 259736 505640 259788 505646
rect 259736 505582 259788 505588
rect 239772 504280 239824 504286
rect 239772 504222 239824 504228
rect 239784 502738 239812 504222
rect 259748 502738 259776 505582
rect 239784 502710 240074 502738
rect 259394 502710 259776 502738
rect 249720 500886 249748 502044
rect 260116 500886 260144 522990
rect 260208 505646 260236 523126
rect 260196 505640 260248 505646
rect 260196 505582 260248 505588
rect 261496 500886 261524 550870
rect 296352 550860 296404 550866
rect 296352 550802 296404 550808
rect 316776 550860 316828 550866
rect 316776 550802 316828 550808
rect 408040 550860 408092 550866
rect 408040 550802 408092 550808
rect 428648 550860 428700 550866
rect 428648 550802 428700 550808
rect 277676 550792 277728 550798
rect 277676 550734 277728 550740
rect 287520 550792 287572 550798
rect 287520 550734 287572 550740
rect 268016 550724 268068 550730
rect 268016 550666 268068 550672
rect 268028 548964 268056 550666
rect 277688 548964 277716 550734
rect 287336 550656 287388 550662
rect 287336 550598 287388 550604
rect 287348 548964 287376 550598
rect 266266 539336 266322 539345
rect 266266 539271 266322 539280
rect 262218 538656 262274 538665
rect 262218 538591 262274 538600
rect 262232 529922 262260 538591
rect 266280 529922 266308 539271
rect 262220 529916 262272 529922
rect 262220 529858 262272 529864
rect 266268 529916 266320 529922
rect 266268 529858 266320 529864
rect 287532 529666 287560 550734
rect 287704 550724 287756 550730
rect 287704 550666 287756 550672
rect 287716 530330 287744 550666
rect 289084 550656 289136 550662
rect 289084 550598 289136 550604
rect 287704 530324 287756 530330
rect 287704 530266 287756 530272
rect 287362 529638 287560 529666
rect 268028 526998 268056 529108
rect 277688 526998 277716 529108
rect 289096 526998 289124 550598
rect 296364 548978 296392 550802
rect 305368 550792 305420 550798
rect 305368 550734 305420 550740
rect 296056 548950 296392 548978
rect 305380 548978 305408 550734
rect 315488 550724 315540 550730
rect 315488 550666 315540 550672
rect 315028 550656 315080 550662
rect 315028 550598 315080 550604
rect 315040 548978 315068 550598
rect 305380 548950 305716 548978
rect 315040 548950 315376 548978
rect 293866 539336 293922 539345
rect 293866 539271 293922 539280
rect 289818 538656 289874 538665
rect 289818 538591 289874 538600
rect 289832 529854 289860 538591
rect 293880 529854 293908 539271
rect 295708 530324 295760 530330
rect 295708 530266 295760 530272
rect 289820 529848 289872 529854
rect 289820 529790 289872 529796
rect 293868 529848 293920 529854
rect 293868 529790 293920 529796
rect 295720 529666 295748 530266
rect 315500 529666 315528 550666
rect 316684 550656 316736 550662
rect 316684 550598 316736 550604
rect 295720 529638 296056 529666
rect 315376 529638 315528 529666
rect 305716 529094 306052 529122
rect 306024 526998 306052 529094
rect 316696 526998 316724 550598
rect 316788 530738 316816 550802
rect 345664 550792 345716 550798
rect 345664 550734 345716 550740
rect 361672 550792 361724 550798
rect 361672 550734 361724 550740
rect 371516 550792 371568 550798
rect 371516 550734 371568 550740
rect 389364 550792 389416 550798
rect 389364 550734 389416 550740
rect 399484 550792 399536 550798
rect 399484 550734 399536 550740
rect 333704 550724 333756 550730
rect 333704 550666 333756 550672
rect 333716 548964 333744 550666
rect 343364 550656 343416 550662
rect 343364 550598 343416 550604
rect 344284 550656 344336 550662
rect 344284 550598 344336 550604
rect 343376 548964 343404 550598
rect 323044 548270 324070 548298
rect 322846 539336 322902 539345
rect 322846 539271 322902 539280
rect 317418 538656 317474 538665
rect 317418 538591 317474 538600
rect 316776 530732 316828 530738
rect 316776 530674 316828 530680
rect 317432 529922 317460 538591
rect 322860 529922 322888 539271
rect 317420 529916 317472 529922
rect 317420 529858 317472 529864
rect 322848 529916 322900 529922
rect 322848 529858 322900 529864
rect 323044 526998 323072 548270
rect 323676 530732 323728 530738
rect 323676 530674 323728 530680
rect 323688 529666 323716 530674
rect 343548 529848 343600 529854
rect 343548 529790 343600 529796
rect 343560 529666 343588 529790
rect 323688 529638 324070 529666
rect 343390 529638 343588 529666
rect 268016 526992 268068 526998
rect 268016 526934 268068 526940
rect 277676 526992 277728 526998
rect 277676 526934 277728 526940
rect 289084 526992 289136 526998
rect 289084 526934 289136 526940
rect 306012 526992 306064 526998
rect 306012 526934 306064 526940
rect 316684 526992 316736 526998
rect 316684 526934 316736 526940
rect 323032 526992 323084 526998
rect 323032 526934 323084 526940
rect 333716 526930 333744 529108
rect 344296 526930 344324 550598
rect 345018 538656 345074 538665
rect 345018 538591 345074 538600
rect 345032 529786 345060 538591
rect 345676 529854 345704 550734
rect 352012 550724 352064 550730
rect 352012 550666 352064 550672
rect 352024 548964 352052 550666
rect 361684 548964 361712 550734
rect 371332 550656 371384 550662
rect 371332 550598 371384 550604
rect 371344 548964 371372 550598
rect 350446 539336 350502 539345
rect 350446 539271 350502 539280
rect 350460 529854 350488 539271
rect 345664 529848 345716 529854
rect 345664 529790 345716 529796
rect 350448 529848 350500 529854
rect 350448 529790 350500 529796
rect 345020 529780 345072 529786
rect 345020 529722 345072 529728
rect 371528 529666 371556 550734
rect 374644 550724 374696 550730
rect 374644 550666 374696 550672
rect 373264 550656 373316 550662
rect 373264 550598 373316 550604
rect 371358 529638 371556 529666
rect 352024 526998 352052 529108
rect 361684 526998 361712 529108
rect 373276 526998 373304 550598
rect 373998 538656 374054 538665
rect 373998 538591 374054 538600
rect 374012 529922 374040 538591
rect 374000 529916 374052 529922
rect 374000 529858 374052 529864
rect 374656 527134 374684 550666
rect 389376 548978 389404 550734
rect 399024 550656 399076 550662
rect 399024 550598 399076 550604
rect 399036 548978 399064 550598
rect 389376 548950 389712 548978
rect 399036 548950 399372 548978
rect 379624 548270 380052 548298
rect 378046 539336 378102 539345
rect 378046 539271 378102 539280
rect 378060 529786 378088 539271
rect 378048 529780 378100 529786
rect 378048 529722 378100 529728
rect 374644 527128 374696 527134
rect 374644 527070 374696 527076
rect 379624 526998 379652 548270
rect 399496 529666 399524 550734
rect 400864 550656 400916 550662
rect 400864 550598 400916 550604
rect 399372 529638 399524 529666
rect 379716 529094 380052 529122
rect 389712 529094 390048 529122
rect 379716 527134 379744 529094
rect 379704 527128 379756 527134
rect 379704 527070 379756 527076
rect 352012 526992 352064 526998
rect 352012 526934 352064 526940
rect 361672 526992 361724 526998
rect 361672 526934 361724 526940
rect 373264 526992 373316 526998
rect 373264 526934 373316 526940
rect 379612 526992 379664 526998
rect 379612 526934 379664 526940
rect 390020 526930 390048 529094
rect 400876 526930 400904 550598
rect 408052 548964 408080 550802
rect 417700 550792 417752 550798
rect 417700 550734 417752 550740
rect 417712 548964 417740 550734
rect 428464 550724 428516 550730
rect 428464 550666 428516 550672
rect 427360 550656 427412 550662
rect 427360 550598 427412 550604
rect 427372 548964 427400 550598
rect 405646 539336 405702 539345
rect 405646 539271 405702 539280
rect 401598 538656 401654 538665
rect 401598 538591 401654 538600
rect 401612 529854 401640 538591
rect 405660 529922 405688 539271
rect 428476 538214 428504 550666
rect 428556 550656 428608 550662
rect 428556 550598 428608 550604
rect 427832 538186 428504 538214
rect 405648 529916 405700 529922
rect 405648 529858 405700 529864
rect 401600 529848 401652 529854
rect 401600 529790 401652 529796
rect 427832 529666 427860 538186
rect 427386 529638 427860 529666
rect 408052 526998 408080 529108
rect 417712 526998 417740 529108
rect 428568 526998 428596 550598
rect 428660 530602 428688 550802
rect 456156 550792 456208 550798
rect 456156 550734 456208 550740
rect 473360 550792 473412 550798
rect 473360 550734 473412 550740
rect 483480 550792 483532 550798
rect 483480 550734 483532 550740
rect 445668 550724 445720 550730
rect 445668 550666 445720 550672
rect 445680 548964 445708 550666
rect 455328 550656 455380 550662
rect 455328 550598 455380 550604
rect 456064 550656 456116 550662
rect 456064 550598 456116 550604
rect 455340 548964 455368 550598
rect 434824 548270 436034 548298
rect 434626 539336 434682 539345
rect 434626 539271 434682 539280
rect 429198 538656 429254 538665
rect 429198 538591 429254 538600
rect 428648 530596 428700 530602
rect 428648 530538 428700 530544
rect 429212 529786 429240 538591
rect 434640 529854 434668 539271
rect 434628 529848 434680 529854
rect 434628 529790 434680 529796
rect 429200 529780 429252 529786
rect 429200 529722 429252 529728
rect 434824 526998 434852 548270
rect 455696 533656 455748 533662
rect 455696 533598 455748 533604
rect 435732 530596 435784 530602
rect 435732 530538 435784 530544
rect 435744 529666 435772 530538
rect 455708 529666 455736 533598
rect 435744 529638 436034 529666
rect 455354 529638 455736 529666
rect 408040 526992 408092 526998
rect 408040 526934 408092 526940
rect 417700 526992 417752 526998
rect 417700 526934 417752 526940
rect 428556 526992 428608 526998
rect 428556 526934 428608 526940
rect 434812 526992 434864 526998
rect 434812 526934 434864 526940
rect 445680 526930 445708 529108
rect 456076 526930 456104 550598
rect 456168 533662 456196 550734
rect 464344 550724 464396 550730
rect 464344 550666 464396 550672
rect 464356 548978 464384 550666
rect 464048 548950 464384 548978
rect 473372 548978 473400 550734
rect 483020 550656 483072 550662
rect 483020 550598 483072 550604
rect 483032 548978 483060 550598
rect 473372 548950 473708 548978
rect 483032 548950 483368 548978
rect 462226 539336 462282 539345
rect 462226 539271 462282 539280
rect 458178 538656 458234 538665
rect 458178 538591 458234 538600
rect 456156 533656 456208 533662
rect 456156 533598 456208 533604
rect 458192 529922 458220 538591
rect 458180 529916 458232 529922
rect 458180 529858 458232 529864
rect 462240 529786 462268 539271
rect 462228 529780 462280 529786
rect 462228 529722 462280 529728
rect 483492 529666 483520 550734
rect 483664 550724 483716 550730
rect 483664 550666 483716 550672
rect 483676 530194 483704 550666
rect 485044 550656 485096 550662
rect 485044 550598 485096 550604
rect 483664 530188 483716 530194
rect 483664 530130 483716 530136
rect 483368 529638 483520 529666
rect 463804 529094 464048 529122
rect 473708 529094 474044 529122
rect 463804 526998 463832 529094
rect 474016 526998 474044 529094
rect 485056 526998 485084 550598
rect 489826 539336 489882 539345
rect 489826 539271 489882 539280
rect 485778 538656 485834 538665
rect 485778 538591 485834 538600
rect 485792 529854 485820 538591
rect 489840 529922 489868 539271
rect 489828 529916 489880 529922
rect 489828 529858 489880 529864
rect 485780 529848 485832 529854
rect 485780 529790 485832 529796
rect 463792 526992 463844 526998
rect 463792 526934 463844 526940
rect 474004 526992 474056 526998
rect 474004 526934 474056 526940
rect 485044 526992 485096 526998
rect 485044 526934 485096 526940
rect 333704 526924 333756 526930
rect 333704 526866 333756 526872
rect 344284 526924 344336 526930
rect 344284 526866 344336 526872
rect 390008 526924 390060 526930
rect 390008 526866 390060 526872
rect 400864 526924 400916 526930
rect 400864 526866 400916 526872
rect 445668 526924 445720 526930
rect 445668 526866 445720 526872
rect 456064 526924 456116 526930
rect 456064 526866 456116 526872
rect 296352 523252 296404 523258
rect 296352 523194 296404 523200
rect 316776 523252 316828 523258
rect 316776 523194 316828 523200
rect 408040 523252 408092 523258
rect 408040 523194 408092 523200
rect 428648 523252 428700 523258
rect 428648 523194 428700 523200
rect 277676 523184 277728 523190
rect 277676 523126 277728 523132
rect 287520 523184 287572 523190
rect 287520 523126 287572 523132
rect 268016 523116 268068 523122
rect 268016 523058 268068 523064
rect 268028 521900 268056 523058
rect 277688 521900 277716 523126
rect 287336 523048 287388 523054
rect 287336 522990 287388 522996
rect 287348 521900 287376 522990
rect 262220 520328 262272 520334
rect 262220 520270 262272 520276
rect 262232 511601 262260 520270
rect 266266 512272 266322 512281
rect 266266 512207 266322 512216
rect 262218 511592 262274 511601
rect 262218 511527 262274 511536
rect 266280 503674 266308 512207
rect 266268 503668 266320 503674
rect 266268 503610 266320 503616
rect 287532 502738 287560 523126
rect 287704 523116 287756 523122
rect 287704 523058 287756 523064
rect 287716 504626 287744 523058
rect 289084 523048 289136 523054
rect 289084 522990 289136 522996
rect 287704 504620 287756 504626
rect 287704 504562 287756 504568
rect 287362 502710 287560 502738
rect 249708 500880 249760 500886
rect 249708 500822 249760 500828
rect 260104 500880 260156 500886
rect 260104 500822 260156 500828
rect 261484 500880 261536 500886
rect 261484 500822 261536 500828
rect 268028 500818 268056 502044
rect 277688 500818 277716 502044
rect 289096 500818 289124 522990
rect 296364 521914 296392 523194
rect 305368 523184 305420 523190
rect 305368 523126 305420 523132
rect 296056 521886 296392 521914
rect 305380 521914 305408 523126
rect 315488 523116 315540 523122
rect 315488 523058 315540 523064
rect 315028 523048 315080 523054
rect 315028 522990 315080 522996
rect 315040 521914 315068 522990
rect 305380 521886 305716 521914
rect 315040 521886 315376 521914
rect 289820 520396 289872 520402
rect 289820 520338 289872 520344
rect 289832 511601 289860 520338
rect 293868 520328 293920 520334
rect 293868 520270 293920 520276
rect 293880 512281 293908 520270
rect 293866 512272 293922 512281
rect 293866 512207 293922 512216
rect 289818 511592 289874 511601
rect 289818 511527 289874 511536
rect 295708 504620 295760 504626
rect 295708 504562 295760 504568
rect 295720 502738 295748 504562
rect 315500 502738 315528 523058
rect 316684 523048 316736 523054
rect 316684 522990 316736 522996
rect 295720 502710 296056 502738
rect 315376 502710 315528 502738
rect 305716 502030 306052 502058
rect 306024 500818 306052 502030
rect 316696 500818 316724 522990
rect 316788 503810 316816 523194
rect 345664 523184 345716 523190
rect 345664 523126 345716 523132
rect 361672 523184 361724 523190
rect 361672 523126 361724 523132
rect 371516 523184 371568 523190
rect 371516 523126 371568 523132
rect 389364 523184 389416 523190
rect 389364 523126 389416 523132
rect 399484 523184 399536 523190
rect 399484 523126 399536 523132
rect 333704 523116 333756 523122
rect 333704 523058 333756 523064
rect 333716 521900 333744 523058
rect 343364 523048 343416 523054
rect 343364 522990 343416 522996
rect 344284 523048 344336 523054
rect 344284 522990 344336 522996
rect 343376 521900 343404 522990
rect 323044 521206 324070 521234
rect 322848 520396 322900 520402
rect 322848 520338 322900 520344
rect 322860 512281 322888 520338
rect 322846 512272 322902 512281
rect 322846 512207 322902 512216
rect 317418 511592 317474 511601
rect 317418 511527 317474 511536
rect 316776 503804 316828 503810
rect 316776 503746 316828 503752
rect 317432 503674 317460 511527
rect 317420 503668 317472 503674
rect 317420 503610 317472 503616
rect 323044 500818 323072 521206
rect 323676 503804 323728 503810
rect 323676 503746 323728 503752
rect 323688 502738 323716 503746
rect 323688 502710 324070 502738
rect 238852 500812 238904 500818
rect 238852 500754 238904 500760
rect 268016 500812 268068 500818
rect 268016 500754 268068 500760
rect 277676 500812 277728 500818
rect 277676 500754 277728 500760
rect 289084 500812 289136 500818
rect 289084 500754 289136 500760
rect 306012 500812 306064 500818
rect 306012 500754 306064 500760
rect 316684 500812 316736 500818
rect 316684 500754 316736 500760
rect 323032 500812 323084 500818
rect 323032 500754 323084 500760
rect 333716 500750 333744 502044
rect 343376 500954 343404 502044
rect 343364 500948 343416 500954
rect 343364 500890 343416 500896
rect 344296 500750 344324 522990
rect 345020 520328 345072 520334
rect 345020 520270 345072 520276
rect 345032 511601 345060 520270
rect 345018 511592 345074 511601
rect 345018 511527 345074 511536
rect 345676 500954 345704 523126
rect 352012 523116 352064 523122
rect 352012 523058 352064 523064
rect 352024 521900 352052 523058
rect 361684 521900 361712 523126
rect 371332 523048 371384 523054
rect 371332 522990 371384 522996
rect 371344 521900 371372 522990
rect 350448 520328 350500 520334
rect 350448 520270 350500 520276
rect 350460 512281 350488 520270
rect 350446 512272 350502 512281
rect 350446 512207 350502 512216
rect 371528 502738 371556 523126
rect 374644 523116 374696 523122
rect 374644 523058 374696 523064
rect 373264 523048 373316 523054
rect 373264 522990 373316 522996
rect 371358 502710 371556 502738
rect 345664 500948 345716 500954
rect 345664 500890 345716 500896
rect 352024 500818 352052 502044
rect 361684 500818 361712 502044
rect 373276 500818 373304 522990
rect 374000 520396 374052 520402
rect 374000 520338 374052 520344
rect 374012 511601 374040 520338
rect 373998 511592 374054 511601
rect 373998 511527 374054 511536
rect 374656 500954 374684 523058
rect 389376 521914 389404 523126
rect 399024 523048 399076 523054
rect 399024 522990 399076 522996
rect 399036 521914 399064 522990
rect 389376 521886 389712 521914
rect 399036 521886 399372 521914
rect 379624 521206 380052 521234
rect 378046 512272 378102 512281
rect 378046 512207 378102 512216
rect 378060 503674 378088 512207
rect 378048 503668 378100 503674
rect 378048 503610 378100 503616
rect 374644 500948 374696 500954
rect 374644 500890 374696 500896
rect 379624 500818 379652 521206
rect 399496 502738 399524 523126
rect 400864 523048 400916 523054
rect 400864 522990 400916 522996
rect 399372 502710 399524 502738
rect 379716 502030 380052 502058
rect 389712 502030 390048 502058
rect 379716 500954 379744 502030
rect 379704 500948 379756 500954
rect 379704 500890 379756 500896
rect 352012 500812 352064 500818
rect 352012 500754 352064 500760
rect 361672 500812 361724 500818
rect 361672 500754 361724 500760
rect 373264 500812 373316 500818
rect 373264 500754 373316 500760
rect 379612 500812 379664 500818
rect 379612 500754 379664 500760
rect 390020 500750 390048 502030
rect 400876 500750 400904 522990
rect 408052 521900 408080 523194
rect 417700 523184 417752 523190
rect 417700 523126 417752 523132
rect 417712 521900 417740 523126
rect 428556 523116 428608 523122
rect 428556 523058 428608 523064
rect 427360 523048 427412 523054
rect 427360 522990 427412 522996
rect 428464 523048 428516 523054
rect 428464 522990 428516 522996
rect 427372 521900 427400 522990
rect 401600 520328 401652 520334
rect 401600 520270 401652 520276
rect 407856 520328 407908 520334
rect 407856 520270 407908 520276
rect 401612 511601 401640 520270
rect 407868 512825 407896 520270
rect 407854 512816 407910 512825
rect 407854 512751 407910 512760
rect 401598 511592 401654 511601
rect 401598 511527 401654 511536
rect 427728 503600 427780 503606
rect 427728 503542 427780 503548
rect 427740 502738 427768 503542
rect 427386 502710 427768 502738
rect 408052 500818 408080 502044
rect 417712 500818 417740 502044
rect 428476 500818 428504 522990
rect 428568 503606 428596 523058
rect 428660 504422 428688 523194
rect 456156 523184 456208 523190
rect 456156 523126 456208 523132
rect 473360 523184 473412 523190
rect 473360 523126 473412 523132
rect 483480 523184 483532 523190
rect 483480 523126 483532 523132
rect 445668 523116 445720 523122
rect 445668 523058 445720 523064
rect 445680 521900 445708 523058
rect 455328 523048 455380 523054
rect 455328 522990 455380 522996
rect 456064 523048 456116 523054
rect 456064 522990 456116 522996
rect 455340 521900 455368 522990
rect 434824 521206 436034 521234
rect 434628 520396 434680 520402
rect 434628 520338 434680 520344
rect 434640 512281 434668 520338
rect 434626 512272 434682 512281
rect 434626 512207 434682 512216
rect 429198 511592 429254 511601
rect 429198 511527 429254 511536
rect 428648 504416 428700 504422
rect 428648 504358 428700 504364
rect 429212 503674 429240 511527
rect 429200 503668 429252 503674
rect 429200 503610 429252 503616
rect 428556 503600 428608 503606
rect 428556 503542 428608 503548
rect 434824 500818 434852 521206
rect 455696 505640 455748 505646
rect 455696 505582 455748 505588
rect 435732 504416 435784 504422
rect 435732 504358 435784 504364
rect 435744 502738 435772 504358
rect 455708 502738 455736 505582
rect 435744 502710 436034 502738
rect 455354 502710 455736 502738
rect 408040 500812 408092 500818
rect 408040 500754 408092 500760
rect 417700 500812 417752 500818
rect 417700 500754 417752 500760
rect 428464 500812 428516 500818
rect 428464 500754 428516 500760
rect 434812 500812 434864 500818
rect 434812 500754 434864 500760
rect 445680 500750 445708 502044
rect 456076 500750 456104 522990
rect 456168 505646 456196 523126
rect 464344 523116 464396 523122
rect 464344 523058 464396 523064
rect 464356 521914 464384 523058
rect 464048 521886 464384 521914
rect 473372 521914 473400 523126
rect 483020 523048 483072 523054
rect 483020 522990 483072 522996
rect 483032 521914 483060 522990
rect 473372 521886 473708 521914
rect 483032 521886 483368 521914
rect 458180 520328 458232 520334
rect 458180 520270 458232 520276
rect 458192 511601 458220 520270
rect 462226 512272 462282 512281
rect 462226 512207 462282 512216
rect 458178 511592 458234 511601
rect 458178 511527 458234 511536
rect 456156 505640 456208 505646
rect 456156 505582 456208 505588
rect 462240 503606 462268 512207
rect 462228 503600 462280 503606
rect 462228 503542 462280 503548
rect 483492 502738 483520 523126
rect 483664 523116 483716 523122
rect 483664 523058 483716 523064
rect 483676 504354 483704 523058
rect 485044 523048 485096 523054
rect 485044 522990 485096 522996
rect 483664 504348 483716 504354
rect 483664 504290 483716 504296
rect 483368 502710 483520 502738
rect 463712 502030 464048 502058
rect 473708 502030 474044 502058
rect 463712 500818 463740 502030
rect 474016 500818 474044 502030
rect 485056 500818 485084 522990
rect 485780 520396 485832 520402
rect 485780 520338 485832 520344
rect 485792 511601 485820 520338
rect 489826 512272 489882 512281
rect 489826 512207 489882 512216
rect 485778 511592 485834 511601
rect 485778 511527 485834 511536
rect 489840 503674 489868 512207
rect 489828 503668 489880 503674
rect 489828 503610 489880 503616
rect 463700 500812 463752 500818
rect 463700 500754 463752 500760
rect 474004 500812 474056 500818
rect 474004 500754 474056 500760
rect 485044 500812 485096 500818
rect 485044 500754 485096 500760
rect 333704 500744 333756 500750
rect 333704 500686 333756 500692
rect 344284 500744 344336 500750
rect 344284 500686 344336 500692
rect 390008 500744 390060 500750
rect 390008 500686 390060 500692
rect 400864 500744 400916 500750
rect 400864 500686 400916 500692
rect 445668 500744 445720 500750
rect 445668 500686 445720 500692
rect 456064 500744 456116 500750
rect 456064 500686 456116 500692
rect 261484 497140 261536 497146
rect 261484 497082 261536 497088
rect 249708 497004 249760 497010
rect 249708 496946 249760 496952
rect 260104 497004 260156 497010
rect 260104 496946 260156 496952
rect 249720 494972 249748 496946
rect 259368 496936 259420 496942
rect 259368 496878 259420 496884
rect 259380 494972 259408 496878
rect 238864 494278 240074 494306
rect 238666 485344 238722 485353
rect 238666 485279 238722 485288
rect 238680 475998 238708 485279
rect 238668 475992 238720 475998
rect 238668 475934 238720 475940
rect 238864 473210 238892 494278
rect 260116 480254 260144 496946
rect 260196 496868 260248 496874
rect 260196 496810 260248 496816
rect 259840 480226 260144 480254
rect 239772 476604 239824 476610
rect 239772 476546 239824 476552
rect 239784 475674 239812 476546
rect 259840 475674 259868 480226
rect 239784 475646 240074 475674
rect 259394 475646 259868 475674
rect 238852 473204 238904 473210
rect 238852 473146 238904 473152
rect 249720 473142 249748 475116
rect 260208 473142 260236 496810
rect 249708 473136 249760 473142
rect 249708 473078 249760 473084
rect 260196 473136 260248 473142
rect 260196 473078 260248 473084
rect 249708 469396 249760 469402
rect 249708 469338 249760 469344
rect 260104 469396 260156 469402
rect 260104 469338 260156 469344
rect 249720 467908 249748 469338
rect 259368 469260 259420 469266
rect 259368 469202 259420 469208
rect 259380 467908 259408 469202
rect 238864 467214 240074 467242
rect 238668 466540 238720 466546
rect 238668 466482 238720 466488
rect 238680 458289 238708 466482
rect 238666 458280 238722 458289
rect 238666 458215 238722 458224
rect 238864 445602 238892 467214
rect 260116 451274 260144 469338
rect 260196 469260 260248 469266
rect 260196 469202 260248 469208
rect 259840 451246 260144 451274
rect 239772 449948 239824 449954
rect 239772 449890 239824 449896
rect 239784 448746 239812 449890
rect 259840 448746 259868 451246
rect 239784 448718 240074 448746
rect 259394 448718 259868 448746
rect 249720 445670 249748 448052
rect 260208 445670 260236 469202
rect 261496 445670 261524 497082
rect 408040 497072 408092 497078
rect 408040 497014 408092 497020
rect 428648 497072 428700 497078
rect 428648 497014 428700 497020
rect 277676 497004 277728 497010
rect 277676 496946 277728 496952
rect 287520 497004 287572 497010
rect 287520 496946 287572 496952
rect 305368 497004 305420 497010
rect 305368 496946 305420 496952
rect 315488 497004 315540 497010
rect 315488 496946 315540 496952
rect 333704 497004 333756 497010
rect 333704 496946 333756 496952
rect 345664 497004 345716 497010
rect 345664 496946 345716 496952
rect 361672 497004 361724 497010
rect 361672 496946 361724 496952
rect 371516 497004 371568 497010
rect 371516 496946 371568 496952
rect 389364 497004 389416 497010
rect 389364 496946 389416 496952
rect 399484 497004 399536 497010
rect 399484 496946 399536 496952
rect 268016 496936 268068 496942
rect 268016 496878 268068 496884
rect 268028 494972 268056 496878
rect 277688 494972 277716 496946
rect 287336 496868 287388 496874
rect 287336 496810 287388 496816
rect 287348 494972 287376 496810
rect 266266 485344 266322 485353
rect 266266 485279 266322 485288
rect 262218 484664 262274 484673
rect 262218 484599 262274 484608
rect 262232 476066 262260 484599
rect 266280 476066 266308 485279
rect 262220 476060 262272 476066
rect 262220 476002 262272 476008
rect 266268 476060 266320 476066
rect 266268 476002 266320 476008
rect 287532 475674 287560 496946
rect 287704 496936 287756 496942
rect 287704 496878 287756 496884
rect 296352 496936 296404 496942
rect 296352 496878 296404 496884
rect 287716 476474 287744 496878
rect 289084 496868 289136 496874
rect 289084 496810 289136 496816
rect 287704 476468 287756 476474
rect 287704 476410 287756 476416
rect 287362 475646 287560 475674
rect 268028 473210 268056 475116
rect 277688 473210 277716 475116
rect 289096 473210 289124 496810
rect 296364 494986 296392 496878
rect 296056 494958 296392 494986
rect 305380 494986 305408 496946
rect 315028 496868 315080 496874
rect 315028 496810 315080 496816
rect 315040 494986 315068 496810
rect 305380 494958 305716 494986
rect 315040 494958 315376 494986
rect 293866 485344 293922 485353
rect 293866 485279 293922 485288
rect 289818 484664 289874 484673
rect 289818 484599 289874 484608
rect 289832 475998 289860 484599
rect 293880 475998 293908 485279
rect 295708 476468 295760 476474
rect 295708 476410 295760 476416
rect 289820 475992 289872 475998
rect 289820 475934 289872 475940
rect 293868 475992 293920 475998
rect 293868 475934 293920 475940
rect 295720 475674 295748 476410
rect 315500 475674 315528 496946
rect 316776 496936 316828 496942
rect 316776 496878 316828 496884
rect 316684 496868 316736 496874
rect 316684 496810 316736 496816
rect 295720 475646 296056 475674
rect 315376 475646 315528 475674
rect 305716 475102 306052 475130
rect 306024 473210 306052 475102
rect 316696 473210 316724 496810
rect 316788 476474 316816 496878
rect 333716 494972 333744 496946
rect 343364 496868 343416 496874
rect 343364 496810 343416 496816
rect 344284 496868 344336 496874
rect 344284 496810 344336 496816
rect 343376 494972 343404 496810
rect 323044 494278 324070 494306
rect 322846 485344 322902 485353
rect 322846 485279 322902 485288
rect 317418 484664 317474 484673
rect 317418 484599 317474 484608
rect 316776 476468 316828 476474
rect 316776 476410 316828 476416
rect 317432 476066 317460 484599
rect 322860 476066 322888 485279
rect 317420 476060 317472 476066
rect 317420 476002 317472 476008
rect 322848 476060 322900 476066
rect 322848 476002 322900 476008
rect 323044 473210 323072 494278
rect 323676 476468 323728 476474
rect 323676 476410 323728 476416
rect 323688 475674 323716 476410
rect 343548 475924 343600 475930
rect 343548 475866 343600 475872
rect 343560 475674 343588 475866
rect 323688 475646 324070 475674
rect 343390 475646 343588 475674
rect 268016 473204 268068 473210
rect 268016 473146 268068 473152
rect 277676 473204 277728 473210
rect 277676 473146 277728 473152
rect 289084 473204 289136 473210
rect 289084 473146 289136 473152
rect 306012 473204 306064 473210
rect 306012 473146 306064 473152
rect 316684 473204 316736 473210
rect 316684 473146 316736 473152
rect 323032 473204 323084 473210
rect 323032 473146 323084 473152
rect 333716 473142 333744 475116
rect 344296 473142 344324 496810
rect 345018 484664 345074 484673
rect 345018 484599 345074 484608
rect 345032 475998 345060 484599
rect 345020 475992 345072 475998
rect 345020 475934 345072 475940
rect 345676 475930 345704 496946
rect 352012 496936 352064 496942
rect 352012 496878 352064 496884
rect 352024 494972 352052 496878
rect 361684 494972 361712 496946
rect 371332 496868 371384 496874
rect 371332 496810 371384 496816
rect 371344 494972 371372 496810
rect 350446 485344 350502 485353
rect 350446 485279 350502 485288
rect 350460 475998 350488 485279
rect 350448 475992 350500 475998
rect 350448 475934 350500 475940
rect 345664 475924 345716 475930
rect 345664 475866 345716 475872
rect 371528 475674 371556 496946
rect 374644 496936 374696 496942
rect 374644 496878 374696 496884
rect 373264 496868 373316 496874
rect 373264 496810 373316 496816
rect 371358 475646 371556 475674
rect 352024 473210 352052 475116
rect 361684 473210 361712 475116
rect 373276 473210 373304 496810
rect 373998 484664 374054 484673
rect 373998 484599 374054 484608
rect 374012 476066 374040 484599
rect 374000 476060 374052 476066
rect 374000 476002 374052 476008
rect 374656 473346 374684 496878
rect 389376 494986 389404 496946
rect 399024 496868 399076 496874
rect 399024 496810 399076 496816
rect 399036 494986 399064 496810
rect 389376 494958 389712 494986
rect 399036 494958 399372 494986
rect 379624 494278 380052 494306
rect 378046 485344 378102 485353
rect 378046 485279 378102 485288
rect 378060 475930 378088 485279
rect 378048 475924 378100 475930
rect 378048 475866 378100 475872
rect 374644 473340 374696 473346
rect 374644 473282 374696 473288
rect 379624 473210 379652 494278
rect 399496 475674 399524 496946
rect 400864 496868 400916 496874
rect 400864 496810 400916 496816
rect 399372 475646 399524 475674
rect 379716 475102 380052 475130
rect 389712 475102 390048 475130
rect 379716 473346 379744 475102
rect 379704 473340 379756 473346
rect 379704 473282 379756 473288
rect 352012 473204 352064 473210
rect 352012 473146 352064 473152
rect 361672 473204 361724 473210
rect 361672 473146 361724 473152
rect 373264 473204 373316 473210
rect 373264 473146 373316 473152
rect 379612 473204 379664 473210
rect 379612 473146 379664 473152
rect 390020 473142 390048 475102
rect 400876 473142 400904 496810
rect 408052 494972 408080 497014
rect 417700 497004 417752 497010
rect 417700 496946 417752 496952
rect 417712 494972 417740 496946
rect 428556 496936 428608 496942
rect 428556 496878 428608 496884
rect 427360 496868 427412 496874
rect 427360 496810 427412 496816
rect 428464 496868 428516 496874
rect 428464 496810 428516 496816
rect 427372 494972 427400 496810
rect 405646 485344 405702 485353
rect 405646 485279 405702 485288
rect 401598 484664 401654 484673
rect 401598 484599 401654 484608
rect 401612 475998 401640 484599
rect 405660 476066 405688 485279
rect 405648 476060 405700 476066
rect 405648 476002 405700 476008
rect 401600 475992 401652 475998
rect 401600 475934 401652 475940
rect 427728 475992 427780 475998
rect 427728 475934 427780 475940
rect 427740 475674 427768 475934
rect 427386 475646 427768 475674
rect 408052 473210 408080 475116
rect 417712 473210 417740 475116
rect 428476 473210 428504 496810
rect 428568 475998 428596 496878
rect 428660 476814 428688 497014
rect 456156 497004 456208 497010
rect 456156 496946 456208 496952
rect 473360 497004 473412 497010
rect 473360 496946 473412 496952
rect 483480 497004 483532 497010
rect 483480 496946 483532 496952
rect 445668 496936 445720 496942
rect 445668 496878 445720 496884
rect 445680 494972 445708 496878
rect 455328 496868 455380 496874
rect 455328 496810 455380 496816
rect 456064 496868 456116 496874
rect 456064 496810 456116 496816
rect 455340 494972 455368 496810
rect 434824 494278 436034 494306
rect 434626 485344 434682 485353
rect 434626 485279 434682 485288
rect 429198 484664 429254 484673
rect 429198 484599 429254 484608
rect 428648 476808 428700 476814
rect 428648 476750 428700 476756
rect 428556 475992 428608 475998
rect 428556 475934 428608 475940
rect 429212 475930 429240 484599
rect 434640 475998 434668 485279
rect 434628 475992 434680 475998
rect 434628 475934 434680 475940
rect 429200 475924 429252 475930
rect 429200 475866 429252 475872
rect 434824 473210 434852 494278
rect 455696 477692 455748 477698
rect 455696 477634 455748 477640
rect 435732 476808 435784 476814
rect 435732 476750 435784 476756
rect 435744 475674 435772 476750
rect 455708 475674 455736 477634
rect 435744 475646 436034 475674
rect 455354 475646 455736 475674
rect 408040 473204 408092 473210
rect 408040 473146 408092 473152
rect 417700 473204 417752 473210
rect 417700 473146 417752 473152
rect 428464 473204 428516 473210
rect 428464 473146 428516 473152
rect 434812 473204 434864 473210
rect 434812 473146 434864 473152
rect 445680 473142 445708 475116
rect 456076 473142 456104 496810
rect 456168 477698 456196 496946
rect 464344 496936 464396 496942
rect 464344 496878 464396 496884
rect 464356 494986 464384 496878
rect 464048 494958 464384 494986
rect 473372 494986 473400 496946
rect 483020 496868 483072 496874
rect 483020 496810 483072 496816
rect 483032 494986 483060 496810
rect 473372 494958 473708 494986
rect 483032 494958 483368 494986
rect 462226 485344 462282 485353
rect 462226 485279 462282 485288
rect 458178 484664 458234 484673
rect 458178 484599 458234 484608
rect 456156 477692 456208 477698
rect 456156 477634 456208 477640
rect 458192 476066 458220 484599
rect 458180 476060 458232 476066
rect 458180 476002 458232 476008
rect 462240 475930 462268 485279
rect 462228 475924 462280 475930
rect 462228 475866 462280 475872
rect 483492 475674 483520 496946
rect 483664 496936 483716 496942
rect 483664 496878 483716 496884
rect 483676 476338 483704 496878
rect 485044 496868 485096 496874
rect 485044 496810 485096 496816
rect 483664 476332 483716 476338
rect 483664 476274 483716 476280
rect 483368 475646 483520 475674
rect 463712 475102 464048 475130
rect 473708 475102 474044 475130
rect 463712 473210 463740 475102
rect 474016 473210 474044 475102
rect 485056 473210 485084 496810
rect 489826 485344 489882 485353
rect 489826 485279 489882 485288
rect 485778 484664 485834 484673
rect 485778 484599 485834 484608
rect 485792 475998 485820 484599
rect 489840 476066 489868 485279
rect 489828 476060 489880 476066
rect 489828 476002 489880 476008
rect 485780 475992 485832 475998
rect 485780 475934 485832 475940
rect 463700 473204 463752 473210
rect 463700 473146 463752 473152
rect 474004 473204 474056 473210
rect 474004 473146 474056 473152
rect 485044 473204 485096 473210
rect 485044 473146 485096 473152
rect 333704 473136 333756 473142
rect 333704 473078 333756 473084
rect 344284 473136 344336 473142
rect 344284 473078 344336 473084
rect 390008 473136 390060 473142
rect 390008 473078 390060 473084
rect 400864 473136 400916 473142
rect 400864 473078 400916 473084
rect 445668 473136 445720 473142
rect 445668 473078 445720 473084
rect 456064 473136 456116 473142
rect 456064 473078 456116 473084
rect 296352 469464 296404 469470
rect 296352 469406 296404 469412
rect 316776 469464 316828 469470
rect 316776 469406 316828 469412
rect 408040 469464 408092 469470
rect 408040 469406 408092 469412
rect 428648 469464 428700 469470
rect 428648 469406 428700 469412
rect 277676 469396 277728 469402
rect 277676 469338 277728 469344
rect 287520 469396 287572 469402
rect 287520 469338 287572 469344
rect 268016 469328 268068 469334
rect 268016 469270 268068 469276
rect 268028 467908 268056 469270
rect 277688 467908 277716 469338
rect 287336 469260 287388 469266
rect 287336 469202 287388 469208
rect 287348 467908 287376 469202
rect 262220 466472 262272 466478
rect 262220 466414 262272 466420
rect 266268 466472 266320 466478
rect 266268 466414 266320 466420
rect 262232 457609 262260 466414
rect 266280 458289 266308 466414
rect 266266 458280 266322 458289
rect 266266 458215 266322 458224
rect 262218 457600 262274 457609
rect 262218 457535 262274 457544
rect 287532 448746 287560 469338
rect 287704 469328 287756 469334
rect 287704 469270 287756 469276
rect 287716 449954 287744 469270
rect 289084 469260 289136 469266
rect 289084 469202 289136 469208
rect 287704 449948 287756 449954
rect 287704 449890 287756 449896
rect 287362 448718 287560 448746
rect 249708 445664 249760 445670
rect 249708 445606 249760 445612
rect 260196 445664 260248 445670
rect 260196 445606 260248 445612
rect 261484 445664 261536 445670
rect 261484 445606 261536 445612
rect 268028 445602 268056 448052
rect 277688 445602 277716 448052
rect 289096 445602 289124 469202
rect 296364 467922 296392 469406
rect 305368 469396 305420 469402
rect 305368 469338 305420 469344
rect 296056 467894 296392 467922
rect 305380 467922 305408 469338
rect 315488 469328 315540 469334
rect 315488 469270 315540 469276
rect 315028 469260 315080 469266
rect 315028 469202 315080 469208
rect 315040 467922 315068 469202
rect 305380 467894 305716 467922
rect 315040 467894 315376 467922
rect 289820 466540 289872 466546
rect 289820 466482 289872 466488
rect 293868 466540 293920 466546
rect 293868 466482 293920 466488
rect 289832 457609 289860 466482
rect 293880 458289 293908 466482
rect 293866 458280 293922 458289
rect 293866 458215 293922 458224
rect 289818 457600 289874 457609
rect 289818 457535 289874 457544
rect 295708 449948 295760 449954
rect 295708 449890 295760 449896
rect 295720 448746 295748 449890
rect 315500 448746 315528 469270
rect 316684 469260 316736 469266
rect 316684 469202 316736 469208
rect 295720 448718 296056 448746
rect 315376 448718 315528 448746
rect 305716 448038 306052 448066
rect 306024 445602 306052 448038
rect 316696 445602 316724 469202
rect 316788 449954 316816 469406
rect 345664 469396 345716 469402
rect 345664 469338 345716 469344
rect 361672 469396 361724 469402
rect 361672 469338 361724 469344
rect 371516 469396 371568 469402
rect 371516 469338 371568 469344
rect 389364 469396 389416 469402
rect 389364 469338 389416 469344
rect 399484 469396 399536 469402
rect 399484 469338 399536 469344
rect 333704 469328 333756 469334
rect 333704 469270 333756 469276
rect 333716 467908 333744 469270
rect 343364 469260 343416 469266
rect 343364 469202 343416 469208
rect 344284 469260 344336 469266
rect 344284 469202 344336 469208
rect 343376 467908 343404 469202
rect 323044 467214 324070 467242
rect 317420 466472 317472 466478
rect 317420 466414 317472 466420
rect 322848 466472 322900 466478
rect 322848 466414 322900 466420
rect 317432 457609 317460 466414
rect 322860 458289 322888 466414
rect 322846 458280 322902 458289
rect 322846 458215 322902 458224
rect 317418 457600 317474 457609
rect 317418 457535 317474 457544
rect 316776 449948 316828 449954
rect 316776 449890 316828 449896
rect 323044 445602 323072 467214
rect 323676 449948 323728 449954
rect 323676 449890 323728 449896
rect 323688 448746 323716 449890
rect 323688 448718 324070 448746
rect 343640 448520 343692 448526
rect 343390 448468 343640 448474
rect 343390 448462 343692 448468
rect 343390 448446 343680 448462
rect 238852 445596 238904 445602
rect 238852 445538 238904 445544
rect 268016 445596 268068 445602
rect 268016 445538 268068 445544
rect 277676 445596 277728 445602
rect 277676 445538 277728 445544
rect 289084 445596 289136 445602
rect 289084 445538 289136 445544
rect 306012 445596 306064 445602
rect 306012 445538 306064 445544
rect 316684 445596 316736 445602
rect 316684 445538 316736 445544
rect 323032 445596 323084 445602
rect 323032 445538 323084 445544
rect 333716 445534 333744 448052
rect 344296 445534 344324 469202
rect 345020 466540 345072 466546
rect 345020 466482 345072 466488
rect 345032 457609 345060 466482
rect 345018 457600 345074 457609
rect 345018 457535 345074 457544
rect 345676 448526 345704 469338
rect 352012 469328 352064 469334
rect 352012 469270 352064 469276
rect 352024 467908 352052 469270
rect 361684 467908 361712 469338
rect 371332 469260 371384 469266
rect 371332 469202 371384 469208
rect 371344 467908 371372 469202
rect 350448 466608 350500 466614
rect 350448 466550 350500 466556
rect 350460 458289 350488 466550
rect 350446 458280 350502 458289
rect 350446 458215 350502 458224
rect 371528 448746 371556 469338
rect 374644 469328 374696 469334
rect 374644 469270 374696 469276
rect 373264 469260 373316 469266
rect 373264 469202 373316 469208
rect 371358 448718 371556 448746
rect 345664 448520 345716 448526
rect 345664 448462 345716 448468
rect 352024 445602 352052 448052
rect 361684 445602 361712 448052
rect 373276 445602 373304 469202
rect 374000 466472 374052 466478
rect 374000 466414 374052 466420
rect 374012 457609 374040 466414
rect 373998 457600 374054 457609
rect 373998 457535 374054 457544
rect 374656 445738 374684 469270
rect 389376 467922 389404 469338
rect 399024 469260 399076 469266
rect 399024 469202 399076 469208
rect 399036 467922 399064 469202
rect 389376 467894 389712 467922
rect 399036 467894 399372 467922
rect 379624 467214 380052 467242
rect 378048 466540 378100 466546
rect 378048 466482 378100 466488
rect 378060 458289 378088 466482
rect 378046 458280 378102 458289
rect 378046 458215 378102 458224
rect 374644 445732 374696 445738
rect 374644 445674 374696 445680
rect 379624 445602 379652 467214
rect 399496 448746 399524 469338
rect 400864 469260 400916 469266
rect 400864 469202 400916 469208
rect 399372 448718 399524 448746
rect 379716 448038 380052 448066
rect 389712 448038 390048 448066
rect 379716 445738 379744 448038
rect 379704 445732 379756 445738
rect 379704 445674 379756 445680
rect 352012 445596 352064 445602
rect 352012 445538 352064 445544
rect 361672 445596 361724 445602
rect 361672 445538 361724 445544
rect 373264 445596 373316 445602
rect 373264 445538 373316 445544
rect 379612 445596 379664 445602
rect 379612 445538 379664 445544
rect 390020 445534 390048 448038
rect 400876 445534 400904 469202
rect 408052 467908 408080 469406
rect 417700 469396 417752 469402
rect 417700 469338 417752 469344
rect 417712 467908 417740 469338
rect 428464 469328 428516 469334
rect 428464 469270 428516 469276
rect 427360 469260 427412 469266
rect 427360 469202 427412 469208
rect 427372 467908 427400 469202
rect 401600 466608 401652 466614
rect 401600 466550 401652 466556
rect 401612 457609 401640 466550
rect 405648 466472 405700 466478
rect 405648 466414 405700 466420
rect 405660 458289 405688 466414
rect 405646 458280 405702 458289
rect 405646 458215 405702 458224
rect 401598 457600 401654 457609
rect 401598 457535 401654 457544
rect 428476 451274 428504 469270
rect 428556 469260 428608 469266
rect 428556 469202 428608 469208
rect 427832 451246 428504 451274
rect 427832 448474 427860 451246
rect 427386 448446 427860 448474
rect 408052 445602 408080 448052
rect 417712 445602 417740 448052
rect 428568 445602 428596 469202
rect 428660 450566 428688 469406
rect 456156 469396 456208 469402
rect 456156 469338 456208 469344
rect 473360 469396 473412 469402
rect 473360 469338 473412 469344
rect 483480 469396 483532 469402
rect 483480 469338 483532 469344
rect 445668 469328 445720 469334
rect 445668 469270 445720 469276
rect 445680 467908 445708 469270
rect 455328 469260 455380 469266
rect 455328 469202 455380 469208
rect 456064 469260 456116 469266
rect 456064 469202 456116 469208
rect 455340 467908 455368 469202
rect 434824 467214 436034 467242
rect 429200 466540 429252 466546
rect 429200 466482 429252 466488
rect 434628 466540 434680 466546
rect 434628 466482 434680 466488
rect 429212 457609 429240 466482
rect 434640 458289 434668 466482
rect 434626 458280 434682 458289
rect 434626 458215 434682 458224
rect 429198 457600 429254 457609
rect 429198 457535 429254 457544
rect 428648 450560 428700 450566
rect 428648 450502 428700 450508
rect 434824 445602 434852 467214
rect 435732 450560 435784 450566
rect 435732 450502 435784 450508
rect 435744 448746 435772 450502
rect 455696 449676 455748 449682
rect 455696 449618 455748 449624
rect 455708 448746 455736 449618
rect 435744 448718 436034 448746
rect 455354 448718 455736 448746
rect 408040 445596 408092 445602
rect 408040 445538 408092 445544
rect 417700 445596 417752 445602
rect 417700 445538 417752 445544
rect 428556 445596 428608 445602
rect 428556 445538 428608 445544
rect 434812 445596 434864 445602
rect 434812 445538 434864 445544
rect 445680 445534 445708 448052
rect 456076 445534 456104 469202
rect 456168 449682 456196 469338
rect 464344 469328 464396 469334
rect 464344 469270 464396 469276
rect 464356 467922 464384 469270
rect 464048 467894 464384 467922
rect 473372 467922 473400 469338
rect 483020 469260 483072 469266
rect 483020 469202 483072 469208
rect 483032 467922 483060 469202
rect 473372 467894 473708 467922
rect 483032 467894 483368 467922
rect 462228 466608 462280 466614
rect 462228 466550 462280 466556
rect 458180 466472 458232 466478
rect 458180 466414 458232 466420
rect 458192 457609 458220 466414
rect 462240 458289 462268 466550
rect 462226 458280 462282 458289
rect 462226 458215 462282 458224
rect 458178 457600 458234 457609
rect 458178 457535 458234 457544
rect 456156 449676 456208 449682
rect 456156 449618 456208 449624
rect 483492 448746 483520 469338
rect 483664 469328 483716 469334
rect 483664 469270 483716 469276
rect 483676 450362 483704 469270
rect 485044 469260 485096 469266
rect 485044 469202 485096 469208
rect 483664 450356 483716 450362
rect 483664 450298 483716 450304
rect 483368 448718 483520 448746
rect 463712 448038 464048 448066
rect 473708 448038 474044 448066
rect 463712 445602 463740 448038
rect 474016 445602 474044 448038
rect 485056 445602 485084 469202
rect 485780 466540 485832 466546
rect 485780 466482 485832 466488
rect 485792 457609 485820 466482
rect 489828 466472 489880 466478
rect 489828 466414 489880 466420
rect 489840 458289 489868 466414
rect 489826 458280 489882 458289
rect 489826 458215 489882 458224
rect 485778 457600 485834 457609
rect 485778 457535 485834 457544
rect 463700 445596 463752 445602
rect 463700 445538 463752 445544
rect 474004 445596 474056 445602
rect 474004 445538 474056 445544
rect 485044 445596 485096 445602
rect 485044 445538 485096 445544
rect 333704 445528 333756 445534
rect 333704 445470 333756 445476
rect 344284 445528 344336 445534
rect 344284 445470 344336 445476
rect 390008 445528 390060 445534
rect 390008 445470 390060 445476
rect 400864 445528 400916 445534
rect 400864 445470 400916 445476
rect 445668 445528 445720 445534
rect 445668 445470 445720 445476
rect 456064 445528 456116 445534
rect 456064 445470 456116 445476
rect 296352 443216 296404 443222
rect 296352 443158 296404 443164
rect 316776 443216 316828 443222
rect 316776 443158 316828 443164
rect 408040 443216 408092 443222
rect 408040 443158 408092 443164
rect 428648 443216 428700 443222
rect 428648 443158 428700 443164
rect 260196 443148 260248 443154
rect 260196 443090 260248 443096
rect 277676 443148 277728 443154
rect 277676 443090 277728 443096
rect 287520 443148 287572 443154
rect 287520 443090 287572 443096
rect 249340 443080 249392 443086
rect 249340 443022 249392 443028
rect 249352 440994 249380 443022
rect 259092 443012 259144 443018
rect 259092 442954 259144 442960
rect 260104 443012 260156 443018
rect 260104 442954 260156 442960
rect 259104 440994 259132 442954
rect 249352 440966 249734 440994
rect 259104 440966 259394 440994
rect 238668 440292 238720 440298
rect 238668 440234 238720 440240
rect 238864 440286 240074 440314
rect 238680 431361 238708 440234
rect 238666 431352 238722 431361
rect 238666 431287 238722 431296
rect 238864 419354 238892 440286
rect 259736 427168 259788 427174
rect 259736 427110 259788 427116
rect 239772 423020 239824 423026
rect 239772 422962 239824 422968
rect 239784 421682 239812 422962
rect 259748 421682 259776 427110
rect 239784 421654 240074 421682
rect 259394 421654 259776 421682
rect 238852 419348 238904 419354
rect 238852 419290 238904 419296
rect 249720 419286 249748 421124
rect 260116 419286 260144 442954
rect 260208 427174 260236 443090
rect 268016 443080 268068 443086
rect 268016 443022 268068 443028
rect 268028 440980 268056 443022
rect 277688 440980 277716 443090
rect 287336 443012 287388 443018
rect 287336 442954 287388 442960
rect 287348 440980 287376 442954
rect 266266 431352 266322 431361
rect 266266 431287 266322 431296
rect 262218 430672 262274 430681
rect 262218 430607 262274 430616
rect 260196 427168 260248 427174
rect 260196 427110 260248 427116
rect 262232 422278 262260 430607
rect 266280 422278 266308 431287
rect 262220 422272 262272 422278
rect 262220 422214 262272 422220
rect 266268 422272 266320 422278
rect 266268 422214 266320 422220
rect 287532 421682 287560 443090
rect 287704 443080 287756 443086
rect 287704 443022 287756 443028
rect 287716 423638 287744 443022
rect 289084 443012 289136 443018
rect 289084 442954 289136 442960
rect 287704 423632 287756 423638
rect 287704 423574 287756 423580
rect 287362 421654 287560 421682
rect 268028 419354 268056 421124
rect 277688 419354 277716 421124
rect 289096 419354 289124 442954
rect 296364 440994 296392 443158
rect 305368 443148 305420 443154
rect 305368 443090 305420 443096
rect 296056 440966 296392 440994
rect 305380 440994 305408 443090
rect 315488 443080 315540 443086
rect 315488 443022 315540 443028
rect 315028 443012 315080 443018
rect 315028 442954 315080 442960
rect 315040 440994 315068 442954
rect 305380 440966 305716 440994
rect 315040 440966 315376 440994
rect 289820 440292 289872 440298
rect 289820 440234 289872 440240
rect 293868 440292 293920 440298
rect 293868 440234 293920 440240
rect 289832 430681 289860 440234
rect 293880 431361 293908 440234
rect 293866 431352 293922 431361
rect 293866 431287 293922 431296
rect 289818 430672 289874 430681
rect 289818 430607 289874 430616
rect 295708 423632 295760 423638
rect 295708 423574 295760 423580
rect 295720 421682 295748 423574
rect 315500 421682 315528 443022
rect 316684 443012 316736 443018
rect 316684 442954 316736 442960
rect 295720 421654 296056 421682
rect 315376 421654 315528 421682
rect 305716 421110 306052 421138
rect 306024 419354 306052 421110
rect 316696 419354 316724 442954
rect 316788 423638 316816 443158
rect 345664 443148 345716 443154
rect 345664 443090 345716 443096
rect 361672 443148 361724 443154
rect 361672 443090 361724 443096
rect 371516 443148 371568 443154
rect 371516 443090 371568 443096
rect 389364 443148 389416 443154
rect 389364 443090 389416 443096
rect 399484 443148 399536 443154
rect 399484 443090 399536 443096
rect 333428 443080 333480 443086
rect 333428 443022 333480 443028
rect 333440 440994 333468 443022
rect 342996 443012 343048 443018
rect 342996 442954 343048 442960
rect 344284 443012 344336 443018
rect 344284 442954 344336 442960
rect 343008 440994 343036 442954
rect 333440 440966 333730 440994
rect 343008 440966 343390 440994
rect 323044 440286 324070 440314
rect 322846 431352 322902 431361
rect 322846 431287 322902 431296
rect 317418 430672 317474 430681
rect 317418 430607 317474 430616
rect 316776 423632 316828 423638
rect 316776 423574 316828 423580
rect 317432 422278 317460 430607
rect 322860 422278 322888 431287
rect 317420 422272 317472 422278
rect 317420 422214 317472 422220
rect 322848 422272 322900 422278
rect 322848 422214 322900 422220
rect 323044 419354 323072 440286
rect 323676 423632 323728 423638
rect 323676 423574 323728 423580
rect 323688 421682 323716 423574
rect 343548 422204 343600 422210
rect 343548 422146 343600 422152
rect 343560 421682 343588 422146
rect 323688 421654 324070 421682
rect 343390 421654 343588 421682
rect 268016 419348 268068 419354
rect 268016 419290 268068 419296
rect 277676 419348 277728 419354
rect 277676 419290 277728 419296
rect 289084 419348 289136 419354
rect 289084 419290 289136 419296
rect 306012 419348 306064 419354
rect 306012 419290 306064 419296
rect 316684 419348 316736 419354
rect 316684 419290 316736 419296
rect 323032 419348 323084 419354
rect 323032 419290 323084 419296
rect 333716 419286 333744 421124
rect 344296 419286 344324 442954
rect 345020 440292 345072 440298
rect 345020 440234 345072 440240
rect 345032 430681 345060 440234
rect 345018 430672 345074 430681
rect 345018 430607 345074 430616
rect 345676 422210 345704 443090
rect 352012 443080 352064 443086
rect 352012 443022 352064 443028
rect 352024 440980 352052 443022
rect 361684 440980 361712 443090
rect 371332 443012 371384 443018
rect 371332 442954 371384 442960
rect 371344 440980 371372 442954
rect 350448 440360 350500 440366
rect 350448 440302 350500 440308
rect 350460 431361 350488 440302
rect 350446 431352 350502 431361
rect 350446 431287 350502 431296
rect 345664 422204 345716 422210
rect 345664 422146 345716 422152
rect 371528 421682 371556 443090
rect 374644 443080 374696 443086
rect 374644 443022 374696 443028
rect 373264 443012 373316 443018
rect 373264 442954 373316 442960
rect 371358 421654 371556 421682
rect 352024 419354 352052 421124
rect 361684 419354 361712 421124
rect 373276 419354 373304 442954
rect 373998 430808 374054 430817
rect 373998 430743 374054 430752
rect 374012 422278 374040 430743
rect 374000 422272 374052 422278
rect 374000 422214 374052 422220
rect 374656 419490 374684 443022
rect 389376 440994 389404 443090
rect 399024 443012 399076 443018
rect 399024 442954 399076 442960
rect 399036 440994 399064 442954
rect 389376 440966 389712 440994
rect 399036 440966 399372 440994
rect 378048 440292 378100 440298
rect 378048 440234 378100 440240
rect 379624 440286 380052 440314
rect 378060 431361 378088 440234
rect 378046 431352 378102 431361
rect 378046 431287 378102 431296
rect 374644 419484 374696 419490
rect 374644 419426 374696 419432
rect 379624 419354 379652 440286
rect 399496 421682 399524 443090
rect 400864 443012 400916 443018
rect 400864 442954 400916 442960
rect 399372 421654 399524 421682
rect 379716 421110 380052 421138
rect 389712 421110 390048 421138
rect 379716 419490 379744 421110
rect 379704 419484 379756 419490
rect 379704 419426 379756 419432
rect 352012 419348 352064 419354
rect 352012 419290 352064 419296
rect 361672 419348 361724 419354
rect 361672 419290 361724 419296
rect 373264 419348 373316 419354
rect 373264 419290 373316 419296
rect 379612 419348 379664 419354
rect 379612 419290 379664 419296
rect 390020 419286 390048 421110
rect 400876 419286 400904 442954
rect 408052 440980 408080 443158
rect 417700 443148 417752 443154
rect 417700 443090 417752 443096
rect 417712 440980 417740 443090
rect 428556 443080 428608 443086
rect 428556 443022 428608 443028
rect 427360 443012 427412 443018
rect 427360 442954 427412 442960
rect 428464 443012 428516 443018
rect 428464 442954 428516 442960
rect 427372 440980 427400 442954
rect 401600 440360 401652 440366
rect 401600 440302 401652 440308
rect 401612 430681 401640 440302
rect 405646 431352 405702 431361
rect 405646 431287 405702 431296
rect 401598 430672 401654 430681
rect 401598 430607 401654 430616
rect 405660 422278 405688 431287
rect 405648 422272 405700 422278
rect 405648 422214 405700 422220
rect 427728 421728 427780 421734
rect 427386 421676 427728 421682
rect 427386 421670 427780 421676
rect 427386 421654 427768 421670
rect 408052 419354 408080 421124
rect 417712 419354 417740 421124
rect 428476 419354 428504 442954
rect 428568 421734 428596 443022
rect 428660 422958 428688 443158
rect 456064 443148 456116 443154
rect 456064 443090 456116 443096
rect 473544 443148 473596 443154
rect 473544 443090 473596 443096
rect 483480 443148 483532 443154
rect 483480 443090 483532 443096
rect 445668 443080 445720 443086
rect 445668 443022 445720 443028
rect 445680 440980 445708 443022
rect 455328 443012 455380 443018
rect 455328 442954 455380 442960
rect 455340 440980 455368 442954
rect 429200 440292 429252 440298
rect 429200 440234 429252 440240
rect 434628 440292 434680 440298
rect 434628 440234 434680 440240
rect 434824 440286 436034 440314
rect 429212 430681 429240 440234
rect 434640 431361 434668 440234
rect 434626 431352 434682 431361
rect 434626 431287 434682 431296
rect 429198 430672 429254 430681
rect 429198 430607 429254 430616
rect 428648 422952 428700 422958
rect 428648 422894 428700 422900
rect 428556 421728 428608 421734
rect 428556 421670 428608 421676
rect 434824 419354 434852 440286
rect 435732 422952 435784 422958
rect 435732 422894 435784 422900
rect 435744 421682 435772 422894
rect 456076 422294 456104 443090
rect 464344 443080 464396 443086
rect 464344 443022 464396 443028
rect 456156 443012 456208 443018
rect 456156 442954 456208 442960
rect 455800 422266 456104 422294
rect 455800 421682 455828 422266
rect 435744 421654 436034 421682
rect 455354 421654 455828 421682
rect 408040 419348 408092 419354
rect 408040 419290 408092 419296
rect 417700 419348 417752 419354
rect 417700 419290 417752 419296
rect 428464 419348 428516 419354
rect 428464 419290 428516 419296
rect 434812 419348 434864 419354
rect 434812 419290 434864 419296
rect 445680 419286 445708 421124
rect 456168 419286 456196 442954
rect 464356 440994 464384 443022
rect 464048 440966 464384 440994
rect 473556 440994 473584 443090
rect 483204 443012 483256 443018
rect 483204 442954 483256 442960
rect 483216 440994 483244 442954
rect 473556 440966 473708 440994
rect 483216 440966 483368 440994
rect 462226 431352 462282 431361
rect 462226 431287 462282 431296
rect 458178 430672 458234 430681
rect 458178 430607 458234 430616
rect 458192 422278 458220 430607
rect 462240 422278 462268 431287
rect 458180 422272 458232 422278
rect 458180 422214 458232 422220
rect 462228 422272 462280 422278
rect 462228 422214 462280 422220
rect 483492 421682 483520 443090
rect 483664 443080 483716 443086
rect 483664 443022 483716 443028
rect 483676 423094 483704 443022
rect 485044 443012 485096 443018
rect 485044 442954 485096 442960
rect 483664 423088 483716 423094
rect 483664 423030 483716 423036
rect 483368 421654 483520 421682
rect 463712 421110 464048 421138
rect 473708 421110 474044 421138
rect 463712 419354 463740 421110
rect 474016 419354 474044 421110
rect 485056 419354 485084 442954
rect 485780 440292 485832 440298
rect 485780 440234 485832 440240
rect 489828 440292 489880 440298
rect 489828 440234 489880 440240
rect 485792 430681 485820 440234
rect 489840 431361 489868 440234
rect 489826 431352 489882 431361
rect 489826 431287 489882 431296
rect 485778 430672 485834 430681
rect 485778 430607 485834 430616
rect 463700 419348 463752 419354
rect 463700 419290 463752 419296
rect 474004 419348 474056 419354
rect 474004 419290 474056 419296
rect 485044 419348 485096 419354
rect 485044 419290 485096 419296
rect 249708 419280 249760 419286
rect 249708 419222 249760 419228
rect 260104 419280 260156 419286
rect 260104 419222 260156 419228
rect 333704 419280 333756 419286
rect 333704 419222 333756 419228
rect 344284 419280 344336 419286
rect 344284 419222 344336 419228
rect 390008 419280 390060 419286
rect 390008 419222 390060 419228
rect 400864 419280 400916 419286
rect 400864 419222 400916 419228
rect 445668 419280 445720 419286
rect 445668 419222 445720 419228
rect 456156 419280 456208 419286
rect 456156 419222 456208 419228
rect 261484 415744 261536 415750
rect 261484 415686 261536 415692
rect 249708 415608 249760 415614
rect 249708 415550 249760 415556
rect 260196 415608 260248 415614
rect 260196 415550 260248 415556
rect 249720 413916 249748 415550
rect 259368 415540 259420 415546
rect 259368 415482 259420 415488
rect 259380 413916 259408 415482
rect 260104 415472 260156 415478
rect 260104 415414 260156 415420
rect 238864 413222 240074 413250
rect 238666 404288 238722 404297
rect 238666 404223 238722 404232
rect 238680 394602 238708 404223
rect 238668 394596 238720 394602
rect 238668 394538 238720 394544
rect 238864 391814 238892 413222
rect 259736 398540 259788 398546
rect 259736 398482 259788 398488
rect 239772 395072 239824 395078
rect 239772 395014 239824 395020
rect 239784 394754 239812 395014
rect 259748 394754 259776 398482
rect 239784 394726 240074 394754
rect 259394 394726 259776 394754
rect 238852 391808 238904 391814
rect 238852 391750 238904 391756
rect 249720 391746 249748 394060
rect 260116 391746 260144 415414
rect 260208 398546 260236 415550
rect 260196 398540 260248 398546
rect 260196 398482 260248 398488
rect 249708 391740 249760 391746
rect 249708 391682 249760 391688
rect 260104 391740 260156 391746
rect 260104 391682 260156 391688
rect 260104 389360 260156 389366
rect 260104 389302 260156 389308
rect 249708 389292 249760 389298
rect 249708 389234 249760 389240
rect 249720 386852 249748 389234
rect 259368 389224 259420 389230
rect 259368 389166 259420 389172
rect 259380 386852 259408 389166
rect 239692 386294 240074 386322
rect 238666 377088 238722 377097
rect 238666 377023 238722 377032
rect 238680 368422 238708 377023
rect 239692 373994 239720 386294
rect 260116 373994 260144 389302
rect 260196 389224 260248 389230
rect 260196 389166 260248 389172
rect 238864 373966 239720 373994
rect 259840 373966 260144 373994
rect 238668 368416 238720 368422
rect 238668 368358 238720 368364
rect 238864 365566 238892 373966
rect 239772 369300 239824 369306
rect 239772 369242 239824 369248
rect 239784 367690 239812 369242
rect 259840 367690 259868 373966
rect 239784 367662 240074 367690
rect 259394 367662 259868 367690
rect 249720 365634 249748 367132
rect 260208 365634 260236 389166
rect 260746 376000 260802 376009
rect 260746 375935 260802 375944
rect 260760 368490 260788 375935
rect 260748 368484 260800 368490
rect 260748 368426 260800 368432
rect 261496 365634 261524 415686
rect 408040 415676 408092 415682
rect 408040 415618 408092 415624
rect 428648 415676 428700 415682
rect 428648 415618 428700 415624
rect 277676 415608 277728 415614
rect 277676 415550 277728 415556
rect 287520 415608 287572 415614
rect 287520 415550 287572 415556
rect 305368 415608 305420 415614
rect 305368 415550 305420 415556
rect 315488 415608 315540 415614
rect 315488 415550 315540 415556
rect 333704 415608 333756 415614
rect 333704 415550 333756 415556
rect 345664 415608 345716 415614
rect 345664 415550 345716 415556
rect 361672 415608 361724 415614
rect 361672 415550 361724 415556
rect 371516 415608 371568 415614
rect 371516 415550 371568 415556
rect 389364 415608 389416 415614
rect 389364 415550 389416 415556
rect 399484 415608 399536 415614
rect 399484 415550 399536 415556
rect 268016 415540 268068 415546
rect 268016 415482 268068 415488
rect 268028 413916 268056 415482
rect 277688 413916 277716 415550
rect 287336 415472 287388 415478
rect 287336 415414 287388 415420
rect 287348 413916 287376 415414
rect 266266 404288 266322 404297
rect 266266 404223 266322 404232
rect 262218 403608 262274 403617
rect 262218 403543 262274 403552
rect 262232 394670 262260 403543
rect 266280 394670 266308 404223
rect 287532 394754 287560 415550
rect 287704 415540 287756 415546
rect 287704 415482 287756 415488
rect 296352 415540 296404 415546
rect 296352 415482 296404 415488
rect 287716 395146 287744 415482
rect 289084 415472 289136 415478
rect 289084 415414 289136 415420
rect 287704 395140 287756 395146
rect 287704 395082 287756 395088
rect 287362 394726 287560 394754
rect 262220 394664 262272 394670
rect 262220 394606 262272 394612
rect 266268 394664 266320 394670
rect 266268 394606 266320 394612
rect 268028 391814 268056 394060
rect 277688 391814 277716 394060
rect 289096 391814 289124 415414
rect 296364 413930 296392 415482
rect 296056 413902 296392 413930
rect 305380 413930 305408 415550
rect 315028 415472 315080 415478
rect 315028 415414 315080 415420
rect 315040 413930 315068 415414
rect 305380 413902 305716 413930
rect 315040 413902 315376 413930
rect 293866 404288 293922 404297
rect 293866 404223 293922 404232
rect 289818 403608 289874 403617
rect 289818 403543 289874 403552
rect 289832 394602 289860 403543
rect 293880 394602 293908 404223
rect 295800 395140 295852 395146
rect 295800 395082 295852 395088
rect 295812 394754 295840 395082
rect 315500 394754 315528 415550
rect 316776 415540 316828 415546
rect 316776 415482 316828 415488
rect 316684 415472 316736 415478
rect 316684 415414 316736 415420
rect 295812 394726 296056 394754
rect 315376 394726 315528 394754
rect 289820 394596 289872 394602
rect 289820 394538 289872 394544
rect 293868 394596 293920 394602
rect 293868 394538 293920 394544
rect 305716 394046 306052 394074
rect 306024 391814 306052 394046
rect 316696 391814 316724 415414
rect 316788 395146 316816 415482
rect 333716 413916 333744 415550
rect 343364 415472 343416 415478
rect 343364 415414 343416 415420
rect 344284 415472 344336 415478
rect 344284 415414 344336 415420
rect 343376 413916 343404 415414
rect 323044 413222 324070 413250
rect 322846 404288 322902 404297
rect 322846 404223 322902 404232
rect 317418 403608 317474 403617
rect 317418 403543 317474 403552
rect 316776 395140 316828 395146
rect 316776 395082 316828 395088
rect 317432 394670 317460 403543
rect 322860 394670 322888 404223
rect 317420 394664 317472 394670
rect 317420 394606 317472 394612
rect 322848 394664 322900 394670
rect 322848 394606 322900 394612
rect 323044 391814 323072 413222
rect 323676 395140 323728 395146
rect 323676 395082 323728 395088
rect 323688 394754 323716 395082
rect 323688 394726 324070 394754
rect 343390 394602 343680 394618
rect 343390 394596 343692 394602
rect 343390 394590 343640 394596
rect 343640 394538 343692 394544
rect 268016 391808 268068 391814
rect 268016 391750 268068 391756
rect 277676 391808 277728 391814
rect 277676 391750 277728 391756
rect 289084 391808 289136 391814
rect 289084 391750 289136 391756
rect 306012 391808 306064 391814
rect 306012 391750 306064 391756
rect 316684 391808 316736 391814
rect 316684 391750 316736 391756
rect 323032 391808 323084 391814
rect 323032 391750 323084 391756
rect 333716 391746 333744 394060
rect 344296 391746 344324 415414
rect 345018 403608 345074 403617
rect 345018 403543 345074 403552
rect 345032 394534 345060 403543
rect 345676 394602 345704 415550
rect 352012 415540 352064 415546
rect 352012 415482 352064 415488
rect 352024 413916 352052 415482
rect 361684 413916 361712 415550
rect 371332 415472 371384 415478
rect 371332 415414 371384 415420
rect 371344 413916 371372 415414
rect 350446 404288 350502 404297
rect 350446 404223 350502 404232
rect 350460 394602 350488 404223
rect 371528 394754 371556 415550
rect 374644 415540 374696 415546
rect 374644 415482 374696 415488
rect 373264 415472 373316 415478
rect 373264 415414 373316 415420
rect 371358 394726 371556 394754
rect 345664 394596 345716 394602
rect 345664 394538 345716 394544
rect 350448 394596 350500 394602
rect 350448 394538 350500 394544
rect 345020 394528 345072 394534
rect 345020 394470 345072 394476
rect 352024 391814 352052 394060
rect 361684 391814 361712 394060
rect 373276 391814 373304 415414
rect 373998 403608 374054 403617
rect 373998 403543 374054 403552
rect 374012 394670 374040 403543
rect 374000 394664 374052 394670
rect 374000 394606 374052 394612
rect 374656 391950 374684 415482
rect 389376 413930 389404 415550
rect 399024 415472 399076 415478
rect 399024 415414 399076 415420
rect 399036 413930 399064 415414
rect 389376 413902 389712 413930
rect 399036 413902 399372 413930
rect 379624 413222 380052 413250
rect 378046 404288 378102 404297
rect 378046 404223 378102 404232
rect 378060 394534 378088 404223
rect 378048 394528 378100 394534
rect 378048 394470 378100 394476
rect 374644 391944 374696 391950
rect 374644 391886 374696 391892
rect 379624 391814 379652 413222
rect 399496 394754 399524 415550
rect 400864 415472 400916 415478
rect 400864 415414 400916 415420
rect 399372 394726 399524 394754
rect 379716 394046 380052 394074
rect 389712 394046 390048 394074
rect 379716 391950 379744 394046
rect 379704 391944 379756 391950
rect 379704 391886 379756 391892
rect 352012 391808 352064 391814
rect 352012 391750 352064 391756
rect 361672 391808 361724 391814
rect 361672 391750 361724 391756
rect 373264 391808 373316 391814
rect 373264 391750 373316 391756
rect 379612 391808 379664 391814
rect 379612 391750 379664 391756
rect 390020 391746 390048 394046
rect 400876 391746 400904 415414
rect 408052 413916 408080 415618
rect 417700 415608 417752 415614
rect 417700 415550 417752 415556
rect 417712 413916 417740 415550
rect 428556 415540 428608 415546
rect 428556 415482 428608 415488
rect 427360 415472 427412 415478
rect 427360 415414 427412 415420
rect 428464 415472 428516 415478
rect 428464 415414 428516 415420
rect 427372 413916 427400 415414
rect 405646 404288 405702 404297
rect 405646 404223 405702 404232
rect 401598 403608 401654 403617
rect 401598 403543 401654 403552
rect 401612 394602 401640 403543
rect 405660 394670 405688 404223
rect 405648 394664 405700 394670
rect 405648 394606 405700 394612
rect 427386 394602 427768 394618
rect 401600 394596 401652 394602
rect 427386 394596 427780 394602
rect 427386 394590 427728 394596
rect 401600 394538 401652 394544
rect 427728 394538 427780 394544
rect 408052 391814 408080 394060
rect 417712 391814 417740 394060
rect 428476 391814 428504 415414
rect 428568 394602 428596 415482
rect 428660 395350 428688 415618
rect 456156 415608 456208 415614
rect 456156 415550 456208 415556
rect 473360 415608 473412 415614
rect 473360 415550 473412 415556
rect 483480 415608 483532 415614
rect 483480 415550 483532 415556
rect 445668 415540 445720 415546
rect 445668 415482 445720 415488
rect 445680 413916 445708 415482
rect 455328 415472 455380 415478
rect 455328 415414 455380 415420
rect 456064 415472 456116 415478
rect 456064 415414 456116 415420
rect 455340 413916 455368 415414
rect 434824 413222 436034 413250
rect 434626 404288 434682 404297
rect 434626 404223 434682 404232
rect 429198 403608 429254 403617
rect 429198 403543 429254 403552
rect 428648 395344 428700 395350
rect 428648 395286 428700 395292
rect 428556 394596 428608 394602
rect 428556 394538 428608 394544
rect 429212 394534 429240 403543
rect 434640 394534 434668 404223
rect 429200 394528 429252 394534
rect 429200 394470 429252 394476
rect 434628 394528 434680 394534
rect 434628 394470 434680 394476
rect 434824 391814 434852 413222
rect 455696 398540 455748 398546
rect 455696 398482 455748 398488
rect 435732 395344 435784 395350
rect 435732 395286 435784 395292
rect 435744 394754 435772 395286
rect 455708 394754 455736 398482
rect 435744 394726 436034 394754
rect 455354 394726 455736 394754
rect 408040 391808 408092 391814
rect 408040 391750 408092 391756
rect 417700 391808 417752 391814
rect 417700 391750 417752 391756
rect 428464 391808 428516 391814
rect 428464 391750 428516 391756
rect 434812 391808 434864 391814
rect 434812 391750 434864 391756
rect 445680 391746 445708 394060
rect 456076 391746 456104 415414
rect 456168 398546 456196 415550
rect 464344 415540 464396 415546
rect 464344 415482 464396 415488
rect 464356 413930 464384 415482
rect 464048 413902 464384 413930
rect 473372 413930 473400 415550
rect 483020 415472 483072 415478
rect 483020 415414 483072 415420
rect 483032 413930 483060 415414
rect 473372 413902 473708 413930
rect 483032 413902 483368 413930
rect 462226 404288 462282 404297
rect 462226 404223 462282 404232
rect 458178 403608 458234 403617
rect 458178 403543 458234 403552
rect 456156 398540 456208 398546
rect 456156 398482 456208 398488
rect 458192 394670 458220 403543
rect 458180 394664 458232 394670
rect 458180 394606 458232 394612
rect 462240 394602 462268 404223
rect 483492 394754 483520 415550
rect 483664 415540 483716 415546
rect 483664 415482 483716 415488
rect 483676 395078 483704 415482
rect 485044 415472 485096 415478
rect 485044 415414 485096 415420
rect 483664 395072 483716 395078
rect 483664 395014 483716 395020
rect 483368 394726 483520 394754
rect 462228 394596 462280 394602
rect 462228 394538 462280 394544
rect 463804 394046 464048 394074
rect 473708 394046 474044 394074
rect 463804 391814 463832 394046
rect 474016 391814 474044 394046
rect 485056 391814 485084 415414
rect 489826 404288 489882 404297
rect 489826 404223 489882 404232
rect 485778 403608 485834 403617
rect 485778 403543 485834 403552
rect 485792 394534 485820 403543
rect 489840 394670 489868 404223
rect 489828 394664 489880 394670
rect 489828 394606 489880 394612
rect 485780 394528 485832 394534
rect 485780 394470 485832 394476
rect 463792 391808 463844 391814
rect 463792 391750 463844 391756
rect 474004 391808 474056 391814
rect 474004 391750 474056 391756
rect 485044 391808 485096 391814
rect 485044 391750 485096 391756
rect 333704 391740 333756 391746
rect 333704 391682 333756 391688
rect 344284 391740 344336 391746
rect 344284 391682 344336 391688
rect 390008 391740 390060 391746
rect 390008 391682 390060 391688
rect 400864 391740 400916 391746
rect 400864 391682 400916 391688
rect 445668 391740 445720 391746
rect 445668 391682 445720 391688
rect 456064 391740 456116 391746
rect 456064 391682 456116 391688
rect 296352 389428 296404 389434
rect 296352 389370 296404 389376
rect 316776 389428 316828 389434
rect 316776 389370 316828 389376
rect 408040 389428 408092 389434
rect 408040 389370 408092 389376
rect 428648 389428 428700 389434
rect 428648 389370 428700 389376
rect 277676 389360 277728 389366
rect 277676 389302 277728 389308
rect 287520 389360 287572 389366
rect 287520 389302 287572 389308
rect 268016 389292 268068 389298
rect 268016 389234 268068 389240
rect 268028 386852 268056 389234
rect 277688 386852 277716 389302
rect 287336 389224 287388 389230
rect 287336 389166 287388 389172
rect 287348 386852 287376 389166
rect 266266 377088 266322 377097
rect 266266 377023 266322 377032
rect 266280 368490 266308 377023
rect 266268 368484 266320 368490
rect 266268 368426 266320 368432
rect 287532 367690 287560 389302
rect 287704 389292 287756 389298
rect 287704 389234 287756 389240
rect 287716 368898 287744 389234
rect 289084 389224 289136 389230
rect 289084 389166 289136 389172
rect 287704 368892 287756 368898
rect 287704 368834 287756 368840
rect 287362 367662 287560 367690
rect 249708 365628 249760 365634
rect 249708 365570 249760 365576
rect 260196 365628 260248 365634
rect 260196 365570 260248 365576
rect 261484 365628 261536 365634
rect 261484 365570 261536 365576
rect 268028 365566 268056 367132
rect 277688 365566 277716 367132
rect 289096 365566 289124 389166
rect 296364 386866 296392 389370
rect 305368 389360 305420 389366
rect 305368 389302 305420 389308
rect 296056 386838 296392 386866
rect 305380 386866 305408 389302
rect 315488 389292 315540 389298
rect 315488 389234 315540 389240
rect 315028 389224 315080 389230
rect 315028 389166 315080 389172
rect 315040 386866 315068 389166
rect 305380 386838 305716 386866
rect 315040 386838 315376 386866
rect 293866 376816 293922 376825
rect 293866 376751 293922 376760
rect 289818 376000 289874 376009
rect 289818 375935 289874 375944
rect 289832 368422 289860 375935
rect 293880 368422 293908 376751
rect 295708 368892 295760 368898
rect 295708 368834 295760 368840
rect 289820 368416 289872 368422
rect 289820 368358 289872 368364
rect 293868 368416 293920 368422
rect 293868 368358 293920 368364
rect 295720 367690 295748 368834
rect 315500 367690 315528 389234
rect 316684 389224 316736 389230
rect 316684 389166 316736 389172
rect 295720 367662 296056 367690
rect 315376 367662 315528 367690
rect 305716 367118 306052 367146
rect 306024 365566 306052 367118
rect 316696 365566 316724 389166
rect 316788 368898 316816 389370
rect 345664 389360 345716 389366
rect 345664 389302 345716 389308
rect 361672 389360 361724 389366
rect 361672 389302 361724 389308
rect 371516 389360 371568 389366
rect 371516 389302 371568 389308
rect 389364 389360 389416 389366
rect 389364 389302 389416 389308
rect 399484 389360 399536 389366
rect 399484 389302 399536 389308
rect 333704 389292 333756 389298
rect 333704 389234 333756 389240
rect 333716 386852 333744 389234
rect 343364 389224 343416 389230
rect 343364 389166 343416 389172
rect 344284 389224 344336 389230
rect 344284 389166 344336 389172
rect 343376 386852 343404 389166
rect 323596 386294 324070 386322
rect 322846 376816 322902 376825
rect 322846 376751 322902 376760
rect 317418 376000 317474 376009
rect 317418 375935 317474 375944
rect 316776 368892 316828 368898
rect 316776 368834 316828 368840
rect 317432 368490 317460 375935
rect 322860 368490 322888 376751
rect 323596 373994 323624 386294
rect 323044 373966 323624 373994
rect 317420 368484 317472 368490
rect 317420 368426 317472 368432
rect 322848 368484 322900 368490
rect 322848 368426 322900 368432
rect 323044 365566 323072 373966
rect 323676 368892 323728 368898
rect 323676 368834 323728 368840
rect 323688 367690 323716 368834
rect 323688 367662 324070 367690
rect 238852 365560 238904 365566
rect 238852 365502 238904 365508
rect 268016 365560 268068 365566
rect 268016 365502 268068 365508
rect 277676 365560 277728 365566
rect 277676 365502 277728 365508
rect 289084 365560 289136 365566
rect 289084 365502 289136 365508
rect 306012 365560 306064 365566
rect 306012 365502 306064 365508
rect 316684 365560 316736 365566
rect 316684 365502 316736 365508
rect 323032 365560 323084 365566
rect 323032 365502 323084 365508
rect 333716 365498 333744 367132
rect 343390 367118 343588 367146
rect 343560 367062 343588 367118
rect 343548 367056 343600 367062
rect 343548 366998 343600 367004
rect 344296 365498 344324 389166
rect 345018 376000 345074 376009
rect 345018 375935 345074 375944
rect 345032 368422 345060 375935
rect 345020 368416 345072 368422
rect 345020 368358 345072 368364
rect 345676 367062 345704 389302
rect 352012 389292 352064 389298
rect 352012 389234 352064 389240
rect 352024 386852 352052 389234
rect 361684 386852 361712 389302
rect 371332 389224 371384 389230
rect 371332 389166 371384 389172
rect 371344 386852 371372 389166
rect 350446 376816 350502 376825
rect 350446 376751 350502 376760
rect 350460 368354 350488 376751
rect 350448 368348 350500 368354
rect 350448 368290 350500 368296
rect 371528 367690 371556 389302
rect 374644 389292 374696 389298
rect 374644 389234 374696 389240
rect 373264 389224 373316 389230
rect 373264 389166 373316 389172
rect 371358 367662 371556 367690
rect 345664 367056 345716 367062
rect 345664 366998 345716 367004
rect 352024 365566 352052 367132
rect 361684 365566 361712 367132
rect 373276 365566 373304 389166
rect 373998 376000 374054 376009
rect 373998 375935 374054 375944
rect 374012 368490 374040 375935
rect 374000 368484 374052 368490
rect 374000 368426 374052 368432
rect 374656 365702 374684 389234
rect 389376 386866 389404 389302
rect 399024 389224 399076 389230
rect 399024 389166 399076 389172
rect 399036 386866 399064 389166
rect 389376 386838 389712 386866
rect 399036 386838 399372 386866
rect 379624 386294 380052 386322
rect 378046 376816 378102 376825
rect 378046 376751 378102 376760
rect 378060 368422 378088 376751
rect 378048 368416 378100 368422
rect 378048 368358 378100 368364
rect 374644 365696 374696 365702
rect 374644 365638 374696 365644
rect 379624 365566 379652 386294
rect 399496 367690 399524 389302
rect 400864 389224 400916 389230
rect 400864 389166 400916 389172
rect 399372 367662 399524 367690
rect 379716 367118 380052 367146
rect 389712 367118 390048 367146
rect 379716 365702 379744 367118
rect 379704 365696 379756 365702
rect 379704 365638 379756 365644
rect 352012 365560 352064 365566
rect 352012 365502 352064 365508
rect 361672 365560 361724 365566
rect 361672 365502 361724 365508
rect 373264 365560 373316 365566
rect 373264 365502 373316 365508
rect 379612 365560 379664 365566
rect 379612 365502 379664 365508
rect 390020 365498 390048 367118
rect 400876 365498 400904 389166
rect 408052 386852 408080 389370
rect 417700 389360 417752 389366
rect 417700 389302 417752 389308
rect 417712 386852 417740 389302
rect 428556 389292 428608 389298
rect 428556 389234 428608 389240
rect 427360 389224 427412 389230
rect 427360 389166 427412 389172
rect 428464 389224 428516 389230
rect 428464 389166 428516 389172
rect 427372 386852 427400 389166
rect 405646 376816 405702 376825
rect 405646 376751 405702 376760
rect 401598 376000 401654 376009
rect 401598 375935 401654 375944
rect 401612 368354 401640 375935
rect 405660 368490 405688 376751
rect 405648 368484 405700 368490
rect 405648 368426 405700 368432
rect 401600 368348 401652 368354
rect 401600 368290 401652 368296
rect 427728 368348 427780 368354
rect 427728 368290 427780 368296
rect 427740 367690 427768 368290
rect 427386 367662 427768 367690
rect 408052 365566 408080 367132
rect 417712 365566 417740 367132
rect 428476 365566 428504 389166
rect 428568 368354 428596 389234
rect 428660 369170 428688 389370
rect 456156 389360 456208 389366
rect 456156 389302 456208 389308
rect 473360 389360 473412 389366
rect 473360 389302 473412 389308
rect 483480 389360 483532 389366
rect 483480 389302 483532 389308
rect 445668 389292 445720 389298
rect 445668 389234 445720 389240
rect 445680 386852 445708 389234
rect 455328 389224 455380 389230
rect 455328 389166 455380 389172
rect 456064 389224 456116 389230
rect 456064 389166 456116 389172
rect 455340 386852 455368 389166
rect 435652 386294 436034 386322
rect 434626 376816 434682 376825
rect 434626 376751 434682 376760
rect 429198 376000 429254 376009
rect 429198 375935 429254 375944
rect 428648 369164 428700 369170
rect 428648 369106 428700 369112
rect 429212 368422 429240 375935
rect 429200 368416 429252 368422
rect 429200 368358 429252 368364
rect 434640 368354 434668 376751
rect 435652 373994 435680 386294
rect 434824 373966 435680 373994
rect 428556 368348 428608 368354
rect 428556 368290 428608 368296
rect 434628 368348 434680 368354
rect 434628 368290 434680 368296
rect 434824 365566 434852 373966
rect 455696 370592 455748 370598
rect 455696 370534 455748 370540
rect 435732 369164 435784 369170
rect 435732 369106 435784 369112
rect 435744 367690 435772 369106
rect 455708 367690 455736 370534
rect 435744 367662 436034 367690
rect 455354 367662 455736 367690
rect 408040 365560 408092 365566
rect 408040 365502 408092 365508
rect 417700 365560 417752 365566
rect 417700 365502 417752 365508
rect 428464 365560 428516 365566
rect 428464 365502 428516 365508
rect 434812 365560 434864 365566
rect 434812 365502 434864 365508
rect 445680 365498 445708 367132
rect 456076 365498 456104 389166
rect 456168 370598 456196 389302
rect 464344 389292 464396 389298
rect 464344 389234 464396 389240
rect 464356 386866 464384 389234
rect 464048 386838 464384 386866
rect 473372 386866 473400 389302
rect 483020 389224 483072 389230
rect 483020 389166 483072 389172
rect 483032 386866 483060 389166
rect 473372 386838 473708 386866
rect 483032 386838 483368 386866
rect 462226 376816 462282 376825
rect 462226 376751 462282 376760
rect 458178 376000 458234 376009
rect 458178 375935 458234 375944
rect 456156 370592 456208 370598
rect 456156 370534 456208 370540
rect 458192 368490 458220 375935
rect 458180 368484 458232 368490
rect 458180 368426 458232 368432
rect 462240 368422 462268 376751
rect 462228 368416 462280 368422
rect 462228 368358 462280 368364
rect 483492 367690 483520 389302
rect 483664 389292 483716 389298
rect 483664 389234 483716 389240
rect 483676 368898 483704 389234
rect 485044 389224 485096 389230
rect 485044 389166 485096 389172
rect 483664 368892 483716 368898
rect 483664 368834 483716 368840
rect 483368 367662 483520 367690
rect 463712 367118 464048 367146
rect 473708 367118 474044 367146
rect 463712 365566 463740 367118
rect 474016 365566 474044 367118
rect 485056 365566 485084 389166
rect 489826 377088 489882 377097
rect 489826 377023 489882 377032
rect 485778 376000 485834 376009
rect 485778 375935 485834 375944
rect 485792 368354 485820 375935
rect 489840 368490 489868 377023
rect 489828 368484 489880 368490
rect 489828 368426 489880 368432
rect 485780 368348 485832 368354
rect 485780 368290 485832 368296
rect 463700 365560 463752 365566
rect 463700 365502 463752 365508
rect 474004 365560 474056 365566
rect 474004 365502 474056 365508
rect 485044 365560 485096 365566
rect 485044 365502 485096 365508
rect 333704 365492 333756 365498
rect 333704 365434 333756 365440
rect 344284 365492 344336 365498
rect 344284 365434 344336 365440
rect 390008 365492 390060 365498
rect 390008 365434 390060 365440
rect 400864 365492 400916 365498
rect 400864 365434 400916 365440
rect 445668 365492 445720 365498
rect 445668 365434 445720 365440
rect 456064 365492 456116 365498
rect 456064 365434 456116 365440
rect 261484 361888 261536 361894
rect 261484 361830 261536 361836
rect 249708 361752 249760 361758
rect 249708 361694 249760 361700
rect 260104 361752 260156 361758
rect 260104 361694 260156 361700
rect 249720 359924 249748 361694
rect 259368 361684 259420 361690
rect 259368 361626 259420 361632
rect 259380 359924 259408 361626
rect 238864 359230 240074 359258
rect 238666 350296 238722 350305
rect 238666 350231 238722 350240
rect 238680 340814 238708 350231
rect 238668 340808 238720 340814
rect 238668 340750 238720 340756
rect 238864 337958 238892 359230
rect 260116 345014 260144 361694
rect 260196 361616 260248 361622
rect 260196 361558 260248 361564
rect 259840 344986 260144 345014
rect 239772 341420 239824 341426
rect 239772 341362 239824 341368
rect 239784 340762 239812 341362
rect 259840 340762 259868 344986
rect 239784 340734 240074 340762
rect 259394 340734 259868 340762
rect 238852 337952 238904 337958
rect 238852 337894 238904 337900
rect 249720 337890 249748 340068
rect 260208 337890 260236 361558
rect 249708 337884 249760 337890
rect 249708 337826 249760 337832
rect 260196 337884 260248 337890
rect 260196 337826 260248 337832
rect 260196 335504 260248 335510
rect 260196 335446 260248 335452
rect 249708 335436 249760 335442
rect 249708 335378 249760 335384
rect 249720 332860 249748 335378
rect 259368 335368 259420 335374
rect 259368 335310 259420 335316
rect 260104 335368 260156 335374
rect 260104 335310 260156 335316
rect 259380 332860 259408 335310
rect 238864 332302 240074 332330
rect 238666 322960 238722 322969
rect 238666 322895 238722 322904
rect 238680 314634 238708 322895
rect 238668 314628 238720 314634
rect 238668 314570 238720 314576
rect 238864 311710 238892 332302
rect 239772 315172 239824 315178
rect 239772 315114 239824 315120
rect 239784 313698 239812 315114
rect 259736 314560 259788 314566
rect 259736 314502 259788 314508
rect 259748 313698 259776 314502
rect 239784 313670 240074 313698
rect 259394 313670 259776 313698
rect 249720 311778 249748 313140
rect 260116 311778 260144 335310
rect 260208 314566 260236 335446
rect 260196 314560 260248 314566
rect 260196 314502 260248 314508
rect 261496 311778 261524 361830
rect 296352 361820 296404 361826
rect 296352 361762 296404 361768
rect 316776 361820 316828 361826
rect 316776 361762 316828 361768
rect 408040 361820 408092 361826
rect 408040 361762 408092 361768
rect 428648 361820 428700 361826
rect 428648 361762 428700 361768
rect 277676 361752 277728 361758
rect 277676 361694 277728 361700
rect 287520 361752 287572 361758
rect 287520 361694 287572 361700
rect 268016 361684 268068 361690
rect 268016 361626 268068 361632
rect 268028 359924 268056 361626
rect 277688 359924 277716 361694
rect 287336 361616 287388 361622
rect 287336 361558 287388 361564
rect 287348 359924 287376 361558
rect 266266 350296 266322 350305
rect 266266 350231 266322 350240
rect 262218 349616 262274 349625
rect 262218 349551 262274 349560
rect 262232 340882 262260 349551
rect 266280 340882 266308 350231
rect 262220 340876 262272 340882
rect 262220 340818 262272 340824
rect 266268 340876 266320 340882
rect 266268 340818 266320 340824
rect 287532 340762 287560 361694
rect 287704 361684 287756 361690
rect 287704 361626 287756 361632
rect 287716 341562 287744 361626
rect 289084 361616 289136 361622
rect 289084 361558 289136 361564
rect 287704 341556 287756 341562
rect 287704 341498 287756 341504
rect 287362 340734 287560 340762
rect 268028 337958 268056 340068
rect 277688 337958 277716 340068
rect 289096 337958 289124 361558
rect 296364 359938 296392 361762
rect 305368 361752 305420 361758
rect 305368 361694 305420 361700
rect 296056 359910 296392 359938
rect 305380 359938 305408 361694
rect 315488 361684 315540 361690
rect 315488 361626 315540 361632
rect 315028 361616 315080 361622
rect 315028 361558 315080 361564
rect 315040 359938 315068 361558
rect 305380 359910 305716 359938
rect 315040 359910 315376 359938
rect 293866 350296 293922 350305
rect 293866 350231 293922 350240
rect 289818 349616 289874 349625
rect 289818 349551 289874 349560
rect 289832 340814 289860 349551
rect 293880 340814 293908 350231
rect 295708 341556 295760 341562
rect 295708 341498 295760 341504
rect 289820 340808 289872 340814
rect 289820 340750 289872 340756
rect 293868 340808 293920 340814
rect 293868 340750 293920 340756
rect 295720 340762 295748 341498
rect 315500 340762 315528 361626
rect 316684 361616 316736 361622
rect 316684 361558 316736 361564
rect 295720 340734 296056 340762
rect 315376 340734 315528 340762
rect 305716 340054 306052 340082
rect 306024 337958 306052 340054
rect 316696 337958 316724 361558
rect 316788 341970 316816 361762
rect 345664 361752 345716 361758
rect 345664 361694 345716 361700
rect 361672 361752 361724 361758
rect 361672 361694 361724 361700
rect 371516 361752 371568 361758
rect 371516 361694 371568 361700
rect 389364 361752 389416 361758
rect 389364 361694 389416 361700
rect 399484 361752 399536 361758
rect 399484 361694 399536 361700
rect 333704 361684 333756 361690
rect 333704 361626 333756 361632
rect 333716 359924 333744 361626
rect 343364 361616 343416 361622
rect 343364 361558 343416 361564
rect 344284 361616 344336 361622
rect 344284 361558 344336 361564
rect 343376 359924 343404 361558
rect 323044 359230 324070 359258
rect 322846 350296 322902 350305
rect 322846 350231 322902 350240
rect 317418 349616 317474 349625
rect 317418 349551 317474 349560
rect 316776 341964 316828 341970
rect 316776 341906 316828 341912
rect 317432 340882 317460 349551
rect 322860 340882 322888 350231
rect 317420 340876 317472 340882
rect 317420 340818 317472 340824
rect 322848 340876 322900 340882
rect 322848 340818 322900 340824
rect 323044 337958 323072 359230
rect 323676 341964 323728 341970
rect 323676 341906 323728 341912
rect 323688 340762 323716 341906
rect 323688 340734 324070 340762
rect 343390 340746 343680 340762
rect 343390 340740 343692 340746
rect 343390 340734 343640 340740
rect 343640 340682 343692 340688
rect 268016 337952 268068 337958
rect 268016 337894 268068 337900
rect 277676 337952 277728 337958
rect 277676 337894 277728 337900
rect 289084 337952 289136 337958
rect 289084 337894 289136 337900
rect 306012 337952 306064 337958
rect 306012 337894 306064 337900
rect 316684 337952 316736 337958
rect 316684 337894 316736 337900
rect 323032 337952 323084 337958
rect 323032 337894 323084 337900
rect 333716 337890 333744 340068
rect 344296 337890 344324 361558
rect 345018 349616 345074 349625
rect 345018 349551 345074 349560
rect 345032 340814 345060 349551
rect 345020 340808 345072 340814
rect 345020 340750 345072 340756
rect 345676 340746 345704 361694
rect 352012 361684 352064 361690
rect 352012 361626 352064 361632
rect 352024 359924 352052 361626
rect 361684 359924 361712 361694
rect 371332 361616 371384 361622
rect 371332 361558 371384 361564
rect 371344 359924 371372 361558
rect 350446 350296 350502 350305
rect 350446 350231 350502 350240
rect 350460 340814 350488 350231
rect 350448 340808 350500 340814
rect 371528 340762 371556 361694
rect 374644 361684 374696 361690
rect 374644 361626 374696 361632
rect 373264 361616 373316 361622
rect 373264 361558 373316 361564
rect 350448 340750 350500 340756
rect 345664 340740 345716 340746
rect 371358 340734 371556 340762
rect 345664 340682 345716 340688
rect 352024 337958 352052 340068
rect 361684 337958 361712 340068
rect 373276 337958 373304 361558
rect 373998 349616 374054 349625
rect 373998 349551 374054 349560
rect 374012 340882 374040 349551
rect 374000 340876 374052 340882
rect 374000 340818 374052 340824
rect 374656 338094 374684 361626
rect 389376 359938 389404 361694
rect 399024 361616 399076 361622
rect 399024 361558 399076 361564
rect 399036 359938 399064 361558
rect 389376 359910 389712 359938
rect 399036 359910 399372 359938
rect 379624 359230 380052 359258
rect 378046 350296 378102 350305
rect 378046 350231 378102 350240
rect 378060 340746 378088 350231
rect 378048 340740 378100 340746
rect 378048 340682 378100 340688
rect 374644 338088 374696 338094
rect 374644 338030 374696 338036
rect 379624 337958 379652 359230
rect 399496 340762 399524 361694
rect 400864 361616 400916 361622
rect 400864 361558 400916 361564
rect 399372 340734 399524 340762
rect 379716 340054 380052 340082
rect 389712 340054 390048 340082
rect 379716 338094 379744 340054
rect 379704 338088 379756 338094
rect 379704 338030 379756 338036
rect 352012 337952 352064 337958
rect 352012 337894 352064 337900
rect 361672 337952 361724 337958
rect 361672 337894 361724 337900
rect 373264 337952 373316 337958
rect 373264 337894 373316 337900
rect 379612 337952 379664 337958
rect 379612 337894 379664 337900
rect 390020 337890 390048 340054
rect 400876 337890 400904 361558
rect 408052 359924 408080 361762
rect 417700 361752 417752 361758
rect 417700 361694 417752 361700
rect 417712 359924 417740 361694
rect 428556 361684 428608 361690
rect 428556 361626 428608 361632
rect 427360 361616 427412 361622
rect 427360 361558 427412 361564
rect 428464 361616 428516 361622
rect 428464 361558 428516 361564
rect 427372 359924 427400 361558
rect 405646 350296 405702 350305
rect 405646 350231 405702 350240
rect 401598 349616 401654 349625
rect 401598 349551 401654 349560
rect 401612 340814 401640 349551
rect 405660 340882 405688 350231
rect 405648 340876 405700 340882
rect 405648 340818 405700 340824
rect 401600 340808 401652 340814
rect 427728 340808 427780 340814
rect 401600 340750 401652 340756
rect 427386 340756 427728 340762
rect 427386 340750 427780 340756
rect 427386 340734 427768 340750
rect 408052 337958 408080 340068
rect 417712 337958 417740 340068
rect 428476 337958 428504 361558
rect 428568 340814 428596 361626
rect 428660 341562 428688 361762
rect 456064 361752 456116 361758
rect 456064 361694 456116 361700
rect 473360 361752 473412 361758
rect 473360 361694 473412 361700
rect 483480 361752 483532 361758
rect 483480 361694 483532 361700
rect 445668 361684 445720 361690
rect 445668 361626 445720 361632
rect 445680 359924 445708 361626
rect 455328 361616 455380 361622
rect 455328 361558 455380 361564
rect 455340 359924 455368 361558
rect 434824 359230 436034 359258
rect 434626 350296 434682 350305
rect 434626 350231 434682 350240
rect 429198 349616 429254 349625
rect 429198 349551 429254 349560
rect 428648 341556 428700 341562
rect 428648 341498 428700 341504
rect 428556 340808 428608 340814
rect 428556 340750 428608 340756
rect 429212 340746 429240 349551
rect 434640 340814 434668 350231
rect 434628 340808 434680 340814
rect 434628 340750 434680 340756
rect 429200 340740 429252 340746
rect 429200 340682 429252 340688
rect 434824 337958 434852 359230
rect 456076 345014 456104 361694
rect 464344 361684 464396 361690
rect 464344 361626 464396 361632
rect 456156 361616 456208 361622
rect 456156 361558 456208 361564
rect 455800 344986 456104 345014
rect 435732 341556 435784 341562
rect 435732 341498 435784 341504
rect 435744 340762 435772 341498
rect 455800 340762 455828 344986
rect 435744 340734 436034 340762
rect 455354 340734 455828 340762
rect 408040 337952 408092 337958
rect 408040 337894 408092 337900
rect 417700 337952 417752 337958
rect 417700 337894 417752 337900
rect 428464 337952 428516 337958
rect 428464 337894 428516 337900
rect 434812 337952 434864 337958
rect 434812 337894 434864 337900
rect 445680 337890 445708 340068
rect 456168 337890 456196 361558
rect 464356 359938 464384 361626
rect 464048 359910 464384 359938
rect 473372 359938 473400 361694
rect 483020 361616 483072 361622
rect 483020 361558 483072 361564
rect 483032 359938 483060 361558
rect 473372 359910 473708 359938
rect 483032 359910 483368 359938
rect 462226 350296 462282 350305
rect 462226 350231 462282 350240
rect 458178 349616 458234 349625
rect 458178 349551 458234 349560
rect 458192 340882 458220 349551
rect 458180 340876 458232 340882
rect 458180 340818 458232 340824
rect 462240 340746 462268 350231
rect 483492 340762 483520 361694
rect 483664 361684 483716 361690
rect 483664 361626 483716 361632
rect 483676 341426 483704 361626
rect 485044 361616 485096 361622
rect 485044 361558 485096 361564
rect 483664 341420 483716 341426
rect 483664 341362 483716 341368
rect 462228 340740 462280 340746
rect 483368 340734 483520 340762
rect 462228 340682 462280 340688
rect 463712 340054 464048 340082
rect 473708 340054 474044 340082
rect 463712 337958 463740 340054
rect 474016 337958 474044 340054
rect 485056 337958 485084 361558
rect 489826 350296 489882 350305
rect 489826 350231 489882 350240
rect 485778 349616 485834 349625
rect 485778 349551 485834 349560
rect 485792 340814 485820 349551
rect 489840 340882 489868 350231
rect 489828 340876 489880 340882
rect 489828 340818 489880 340824
rect 485780 340808 485832 340814
rect 485780 340750 485832 340756
rect 463700 337952 463752 337958
rect 463700 337894 463752 337900
rect 474004 337952 474056 337958
rect 474004 337894 474056 337900
rect 485044 337952 485096 337958
rect 485044 337894 485096 337900
rect 333704 337884 333756 337890
rect 333704 337826 333756 337832
rect 344284 337884 344336 337890
rect 344284 337826 344336 337832
rect 390008 337884 390060 337890
rect 390008 337826 390060 337832
rect 400864 337884 400916 337890
rect 400864 337826 400916 337832
rect 445668 337884 445720 337890
rect 445668 337826 445720 337832
rect 456156 337884 456208 337890
rect 456156 337826 456208 337832
rect 296352 335572 296404 335578
rect 296352 335514 296404 335520
rect 316776 335572 316828 335578
rect 316776 335514 316828 335520
rect 408040 335572 408092 335578
rect 408040 335514 408092 335520
rect 428648 335572 428700 335578
rect 428648 335514 428700 335520
rect 277676 335504 277728 335510
rect 277676 335446 277728 335452
rect 287520 335504 287572 335510
rect 287520 335446 287572 335452
rect 268016 335436 268068 335442
rect 268016 335378 268068 335384
rect 268028 332860 268056 335378
rect 277688 332860 277716 335446
rect 287336 335368 287388 335374
rect 287336 335310 287388 335316
rect 287348 332860 287376 335310
rect 262220 331288 262272 331294
rect 262220 331230 262272 331236
rect 266268 331288 266320 331294
rect 266268 331230 266320 331236
rect 262232 322833 262260 331230
rect 266280 323921 266308 331230
rect 266266 323912 266322 323921
rect 266266 323847 266322 323856
rect 262218 322824 262274 322833
rect 262218 322759 262274 322768
rect 287532 313698 287560 335446
rect 287704 335436 287756 335442
rect 287704 335378 287756 335384
rect 287716 314702 287744 335378
rect 289084 335368 289136 335374
rect 289084 335310 289136 335316
rect 287704 314696 287756 314702
rect 287704 314638 287756 314644
rect 287362 313670 287560 313698
rect 249708 311772 249760 311778
rect 249708 311714 249760 311720
rect 260104 311772 260156 311778
rect 260104 311714 260156 311720
rect 261484 311772 261536 311778
rect 261484 311714 261536 311720
rect 268028 311710 268056 313140
rect 277688 311710 277716 313140
rect 289096 311710 289124 335310
rect 296364 332874 296392 335514
rect 305368 335504 305420 335510
rect 305368 335446 305420 335452
rect 296056 332846 296392 332874
rect 305380 332874 305408 335446
rect 315488 335436 315540 335442
rect 315488 335378 315540 335384
rect 315028 335368 315080 335374
rect 315028 335310 315080 335316
rect 315040 332874 315068 335310
rect 305380 332846 305716 332874
rect 315040 332846 315376 332874
rect 293866 322960 293922 322969
rect 293866 322895 293922 322904
rect 289818 322008 289874 322017
rect 289818 321943 289874 321952
rect 289832 314634 289860 321943
rect 293880 314634 293908 322895
rect 295708 314696 295760 314702
rect 295708 314638 295760 314644
rect 289820 314628 289872 314634
rect 289820 314570 289872 314576
rect 293868 314628 293920 314634
rect 293868 314570 293920 314576
rect 295720 313698 295748 314638
rect 315500 313698 315528 335378
rect 316684 335368 316736 335374
rect 316684 335310 316736 335316
rect 295720 313670 296056 313698
rect 315376 313670 315528 313698
rect 305716 313126 306052 313154
rect 306024 311710 306052 313126
rect 316696 311710 316724 335310
rect 316788 314702 316816 335514
rect 345664 335504 345716 335510
rect 345664 335446 345716 335452
rect 361672 335504 361724 335510
rect 361672 335446 361724 335452
rect 371516 335504 371568 335510
rect 371516 335446 371568 335452
rect 389364 335504 389416 335510
rect 389364 335446 389416 335452
rect 399484 335504 399536 335510
rect 399484 335446 399536 335452
rect 333704 335436 333756 335442
rect 333704 335378 333756 335384
rect 333716 332860 333744 335378
rect 343364 335368 343416 335374
rect 343364 335310 343416 335316
rect 344284 335368 344336 335374
rect 344284 335310 344336 335316
rect 343376 332860 343404 335310
rect 323044 332302 324070 332330
rect 317420 331288 317472 331294
rect 317420 331230 317472 331236
rect 317432 322833 317460 331230
rect 322846 322960 322902 322969
rect 322846 322895 322902 322904
rect 317418 322824 317474 322833
rect 317418 322759 317474 322768
rect 316776 314696 316828 314702
rect 316776 314638 316828 314644
rect 322860 314566 322888 322895
rect 322848 314560 322900 314566
rect 322848 314502 322900 314508
rect 323044 311710 323072 332302
rect 323676 314696 323728 314702
rect 323676 314638 323728 314644
rect 323688 313698 323716 314638
rect 343548 314492 343600 314498
rect 343548 314434 343600 314440
rect 343560 313698 343588 314434
rect 323688 313670 324070 313698
rect 343390 313670 343588 313698
rect 238852 311704 238904 311710
rect 238852 311646 238904 311652
rect 268016 311704 268068 311710
rect 268016 311646 268068 311652
rect 277676 311704 277728 311710
rect 277676 311646 277728 311652
rect 289084 311704 289136 311710
rect 289084 311646 289136 311652
rect 306012 311704 306064 311710
rect 306012 311646 306064 311652
rect 316684 311704 316736 311710
rect 316684 311646 316736 311652
rect 323032 311704 323084 311710
rect 323032 311646 323084 311652
rect 333716 311642 333744 313140
rect 344296 311642 344324 335310
rect 345018 322008 345074 322017
rect 345018 321943 345074 321952
rect 345032 314634 345060 321943
rect 345020 314628 345072 314634
rect 345020 314570 345072 314576
rect 345676 314498 345704 335446
rect 352012 335436 352064 335442
rect 352012 335378 352064 335384
rect 352024 332860 352052 335378
rect 361684 332860 361712 335446
rect 371332 335368 371384 335374
rect 371332 335310 371384 335316
rect 371344 332860 371372 335310
rect 350446 322960 350502 322969
rect 350446 322895 350502 322904
rect 350460 314634 350488 322895
rect 350448 314628 350500 314634
rect 350448 314570 350500 314576
rect 345664 314492 345716 314498
rect 345664 314434 345716 314440
rect 371528 313698 371556 335446
rect 374644 335436 374696 335442
rect 374644 335378 374696 335384
rect 373264 335368 373316 335374
rect 373264 335310 373316 335316
rect 371358 313670 371556 313698
rect 352024 311710 352052 313140
rect 361684 311710 361712 313140
rect 373276 311710 373304 335310
rect 373998 322008 374054 322017
rect 373998 321943 374054 321952
rect 374012 314566 374040 321943
rect 374000 314560 374052 314566
rect 374000 314502 374052 314508
rect 374656 311846 374684 335378
rect 389376 332874 389404 335446
rect 399024 335368 399076 335374
rect 399024 335310 399076 335316
rect 399036 332874 399064 335310
rect 389376 332846 389712 332874
rect 399036 332846 399372 332874
rect 379624 332302 380052 332330
rect 378046 322960 378102 322969
rect 378046 322895 378102 322904
rect 378060 314566 378088 322895
rect 378048 314560 378100 314566
rect 378048 314502 378100 314508
rect 374644 311840 374696 311846
rect 374644 311782 374696 311788
rect 379624 311710 379652 332302
rect 399496 313698 399524 335446
rect 400864 335368 400916 335374
rect 400864 335310 400916 335316
rect 399372 313670 399524 313698
rect 379716 313126 380052 313154
rect 389712 313126 390048 313154
rect 379716 311846 379744 313126
rect 379704 311840 379756 311846
rect 379704 311782 379756 311788
rect 352012 311704 352064 311710
rect 352012 311646 352064 311652
rect 361672 311704 361724 311710
rect 361672 311646 361724 311652
rect 373264 311704 373316 311710
rect 373264 311646 373316 311652
rect 379612 311704 379664 311710
rect 379612 311646 379664 311652
rect 390020 311642 390048 313126
rect 400876 311642 400904 335310
rect 408052 332860 408080 335514
rect 417700 335504 417752 335510
rect 417700 335446 417752 335452
rect 417712 332860 417740 335446
rect 428556 335436 428608 335442
rect 428556 335378 428608 335384
rect 427360 335368 427412 335374
rect 427360 335310 427412 335316
rect 428464 335368 428516 335374
rect 428464 335310 428516 335316
rect 427372 332860 427400 335310
rect 405648 331288 405700 331294
rect 405648 331230 405700 331236
rect 405660 323921 405688 331230
rect 405646 323912 405702 323921
rect 405646 323847 405702 323856
rect 401598 322008 401654 322017
rect 401598 321943 401654 321952
rect 401612 314634 401640 321943
rect 401600 314628 401652 314634
rect 401600 314570 401652 314576
rect 427728 314628 427780 314634
rect 427728 314570 427780 314576
rect 427740 313698 427768 314570
rect 427386 313670 427768 313698
rect 408052 311710 408080 313140
rect 417712 311710 417740 313140
rect 428476 311710 428504 335310
rect 428568 314634 428596 335378
rect 428660 315314 428688 335514
rect 456156 335504 456208 335510
rect 456156 335446 456208 335452
rect 473544 335504 473596 335510
rect 473544 335446 473596 335452
rect 483480 335504 483532 335510
rect 483480 335446 483532 335452
rect 445668 335436 445720 335442
rect 445668 335378 445720 335384
rect 445680 332860 445708 335378
rect 455328 335368 455380 335374
rect 455328 335310 455380 335316
rect 456064 335368 456116 335374
rect 456064 335310 456116 335316
rect 455340 332860 455368 335310
rect 434824 332302 436034 332330
rect 434626 322960 434682 322969
rect 434626 322895 434682 322904
rect 429198 322008 429254 322017
rect 429198 321943 429254 321952
rect 428648 315308 428700 315314
rect 428648 315250 428700 315256
rect 428556 314628 428608 314634
rect 428556 314570 428608 314576
rect 429212 314566 429240 321943
rect 434640 314634 434668 322895
rect 434628 314628 434680 314634
rect 434628 314570 434680 314576
rect 429200 314560 429252 314566
rect 429200 314502 429252 314508
rect 434824 311710 434852 332302
rect 435732 315308 435784 315314
rect 435732 315250 435784 315256
rect 435744 313698 435772 315250
rect 455696 314560 455748 314566
rect 455696 314502 455748 314508
rect 455708 313698 455736 314502
rect 435744 313670 436034 313698
rect 455354 313670 455736 313698
rect 408040 311704 408092 311710
rect 408040 311646 408092 311652
rect 417700 311704 417752 311710
rect 417700 311646 417752 311652
rect 428464 311704 428516 311710
rect 428464 311646 428516 311652
rect 434812 311704 434864 311710
rect 434812 311646 434864 311652
rect 445680 311642 445708 313140
rect 456076 311642 456104 335310
rect 456168 314566 456196 335446
rect 464344 335436 464396 335442
rect 464344 335378 464396 335384
rect 464356 332874 464384 335378
rect 464048 332846 464384 332874
rect 473556 332874 473584 335446
rect 483204 335368 483256 335374
rect 483204 335310 483256 335316
rect 483216 332874 483244 335310
rect 473556 332846 473708 332874
rect 483216 332846 483368 332874
rect 458180 331288 458232 331294
rect 458180 331230 458232 331236
rect 462228 331288 462280 331294
rect 462228 331230 462280 331236
rect 458192 322833 458220 331230
rect 462240 323921 462268 331230
rect 462226 323912 462282 323921
rect 462226 323847 462282 323856
rect 458178 322824 458234 322833
rect 458178 322759 458234 322768
rect 456156 314560 456208 314566
rect 456156 314502 456208 314508
rect 483492 313698 483520 335446
rect 483664 335436 483716 335442
rect 483664 335378 483716 335384
rect 483676 315994 483704 335378
rect 485044 335368 485096 335374
rect 485044 335310 485096 335316
rect 483664 315988 483716 315994
rect 483664 315930 483716 315936
rect 483368 313670 483520 313698
rect 463712 313126 464048 313154
rect 473708 313126 474044 313154
rect 463712 311710 463740 313126
rect 474016 311710 474044 313126
rect 485056 311710 485084 335310
rect 489826 322960 489882 322969
rect 489826 322895 489882 322904
rect 485778 322008 485834 322017
rect 485778 321943 485834 321952
rect 485792 314634 485820 321943
rect 489840 314634 489868 322895
rect 485780 314628 485832 314634
rect 485780 314570 485832 314576
rect 489828 314628 489880 314634
rect 489828 314570 489880 314576
rect 463700 311704 463752 311710
rect 463700 311646 463752 311652
rect 474004 311704 474056 311710
rect 474004 311646 474056 311652
rect 485044 311704 485096 311710
rect 485044 311646 485096 311652
rect 333704 311636 333756 311642
rect 333704 311578 333756 311584
rect 344284 311636 344336 311642
rect 344284 311578 344336 311584
rect 390008 311636 390060 311642
rect 390008 311578 390060 311584
rect 400864 311636 400916 311642
rect 400864 311578 400916 311584
rect 445668 311636 445720 311642
rect 445668 311578 445720 311584
rect 456064 311636 456116 311642
rect 456064 311578 456116 311584
rect 261484 308100 261536 308106
rect 261484 308042 261536 308048
rect 249708 307964 249760 307970
rect 249708 307906 249760 307912
rect 260196 307964 260248 307970
rect 260196 307906 260248 307912
rect 249720 305932 249748 307906
rect 259368 307896 259420 307902
rect 259368 307838 259420 307844
rect 259380 305932 259408 307838
rect 260104 307828 260156 307834
rect 260104 307770 260156 307776
rect 238864 305238 240074 305266
rect 238666 296304 238722 296313
rect 238666 296239 238722 296248
rect 238680 286958 238708 296239
rect 238668 286952 238720 286958
rect 238668 286894 238720 286900
rect 238864 284170 238892 305238
rect 259736 291916 259788 291922
rect 259736 291858 259788 291864
rect 239772 287972 239824 287978
rect 239772 287914 239824 287920
rect 239784 286770 239812 287914
rect 259748 286770 259776 291858
rect 239784 286742 240074 286770
rect 259394 286742 259776 286770
rect 238852 284164 238904 284170
rect 238852 284106 238904 284112
rect 249720 284102 249748 286076
rect 260116 284102 260144 307770
rect 260208 291922 260236 307906
rect 260196 291916 260248 291922
rect 260196 291858 260248 291864
rect 249708 284096 249760 284102
rect 249708 284038 249760 284044
rect 260104 284096 260156 284102
rect 260104 284038 260156 284044
rect 260104 280356 260156 280362
rect 260104 280298 260156 280304
rect 249708 280288 249760 280294
rect 249708 280230 249760 280236
rect 249720 278868 249748 280230
rect 259368 280220 259420 280226
rect 259368 280162 259420 280168
rect 259380 278868 259408 280162
rect 238864 278310 240074 278338
rect 238668 277500 238720 277506
rect 238668 277442 238720 277448
rect 238680 269249 238708 277442
rect 238666 269240 238722 269249
rect 238666 269175 238722 269184
rect 238864 256562 238892 278310
rect 260116 267734 260144 280298
rect 260196 280220 260248 280226
rect 260196 280162 260248 280168
rect 259840 267706 260144 267734
rect 239772 262200 239824 262206
rect 239772 262142 239824 262148
rect 239784 259706 239812 262142
rect 259840 259706 259868 267706
rect 239784 259678 240074 259706
rect 259394 259678 259868 259706
rect 249720 256630 249748 259148
rect 260208 256630 260236 280162
rect 261496 256630 261524 308042
rect 296352 308032 296404 308038
rect 296352 307974 296404 307980
rect 316776 308032 316828 308038
rect 316776 307974 316828 307980
rect 408040 308032 408092 308038
rect 408040 307974 408092 307980
rect 428648 308032 428700 308038
rect 428648 307974 428700 307980
rect 277676 307964 277728 307970
rect 277676 307906 277728 307912
rect 287520 307964 287572 307970
rect 287520 307906 287572 307912
rect 268016 307896 268068 307902
rect 268016 307838 268068 307844
rect 268028 305932 268056 307838
rect 277688 305932 277716 307906
rect 287336 307828 287388 307834
rect 287336 307770 287388 307776
rect 287348 305932 287376 307770
rect 266266 296304 266322 296313
rect 266266 296239 266322 296248
rect 262218 295624 262274 295633
rect 262218 295559 262274 295568
rect 262232 287026 262260 295559
rect 266280 287026 266308 296239
rect 262220 287020 262272 287026
rect 262220 286962 262272 286968
rect 266268 287020 266320 287026
rect 266268 286962 266320 286968
rect 287532 286770 287560 307906
rect 287704 307896 287756 307902
rect 287704 307838 287756 307844
rect 287716 288386 287744 307838
rect 289084 307828 289136 307834
rect 289084 307770 289136 307776
rect 287704 288380 287756 288386
rect 287704 288322 287756 288328
rect 287362 286742 287560 286770
rect 268028 284170 268056 286076
rect 277688 284170 277716 286076
rect 289096 284170 289124 307770
rect 296364 305946 296392 307974
rect 305368 307964 305420 307970
rect 305368 307906 305420 307912
rect 296056 305918 296392 305946
rect 305380 305946 305408 307906
rect 315488 307896 315540 307902
rect 315488 307838 315540 307844
rect 315028 307828 315080 307834
rect 315028 307770 315080 307776
rect 315040 305946 315068 307770
rect 305380 305918 305716 305946
rect 315040 305918 315376 305946
rect 293866 296304 293922 296313
rect 293866 296239 293922 296248
rect 289818 295624 289874 295633
rect 289818 295559 289874 295568
rect 289832 286958 289860 295559
rect 293880 286958 293908 296239
rect 295708 288380 295760 288386
rect 295708 288322 295760 288328
rect 289820 286952 289872 286958
rect 289820 286894 289872 286900
rect 293868 286952 293920 286958
rect 293868 286894 293920 286900
rect 295720 286770 295748 288322
rect 315500 286770 315528 307838
rect 316684 307828 316736 307834
rect 316684 307770 316736 307776
rect 295720 286742 296056 286770
rect 315376 286742 315528 286770
rect 305716 286062 306052 286090
rect 306024 284170 306052 286062
rect 316696 284170 316724 307770
rect 316788 288386 316816 307974
rect 345664 307964 345716 307970
rect 345664 307906 345716 307912
rect 361672 307964 361724 307970
rect 361672 307906 361724 307912
rect 371516 307964 371568 307970
rect 371516 307906 371568 307912
rect 389364 307964 389416 307970
rect 389364 307906 389416 307912
rect 399484 307964 399536 307970
rect 399484 307906 399536 307912
rect 333704 307896 333756 307902
rect 333704 307838 333756 307844
rect 333716 305932 333744 307838
rect 343364 307828 343416 307834
rect 343364 307770 343416 307776
rect 344284 307828 344336 307834
rect 344284 307770 344336 307776
rect 343376 305932 343404 307770
rect 323044 305238 324070 305266
rect 322846 296304 322902 296313
rect 322846 296239 322902 296248
rect 317418 295624 317474 295633
rect 317418 295559 317474 295568
rect 316776 288380 316828 288386
rect 316776 288322 316828 288328
rect 317432 287026 317460 295559
rect 322860 287026 322888 296239
rect 317420 287020 317472 287026
rect 317420 286962 317472 286968
rect 322848 287020 322900 287026
rect 322848 286962 322900 286968
rect 323044 284170 323072 305238
rect 323676 288380 323728 288386
rect 323676 288322 323728 288328
rect 323688 286770 323716 288322
rect 343548 286952 343600 286958
rect 343548 286894 343600 286900
rect 343560 286770 343588 286894
rect 323688 286742 324070 286770
rect 343390 286742 343588 286770
rect 268016 284164 268068 284170
rect 268016 284106 268068 284112
rect 277676 284164 277728 284170
rect 277676 284106 277728 284112
rect 289084 284164 289136 284170
rect 289084 284106 289136 284112
rect 306012 284164 306064 284170
rect 306012 284106 306064 284112
rect 316684 284164 316736 284170
rect 316684 284106 316736 284112
rect 323032 284164 323084 284170
rect 323032 284106 323084 284112
rect 333716 284102 333744 286076
rect 344296 284102 344324 307770
rect 345018 295624 345074 295633
rect 345018 295559 345074 295568
rect 345032 286890 345060 295559
rect 345676 286958 345704 307906
rect 352012 307896 352064 307902
rect 352012 307838 352064 307844
rect 352024 305932 352052 307838
rect 361684 305932 361712 307906
rect 371332 307828 371384 307834
rect 371332 307770 371384 307776
rect 371344 305932 371372 307770
rect 350446 296304 350502 296313
rect 350446 296239 350502 296248
rect 350460 286958 350488 296239
rect 345664 286952 345716 286958
rect 345664 286894 345716 286900
rect 350448 286952 350500 286958
rect 350448 286894 350500 286900
rect 345020 286884 345072 286890
rect 345020 286826 345072 286832
rect 371528 286770 371556 307906
rect 374644 307896 374696 307902
rect 374644 307838 374696 307844
rect 373264 307828 373316 307834
rect 373264 307770 373316 307776
rect 371358 286742 371556 286770
rect 352024 284170 352052 286076
rect 361684 284170 361712 286076
rect 373276 284170 373304 307770
rect 373998 295624 374054 295633
rect 373998 295559 374054 295568
rect 374012 287026 374040 295559
rect 374000 287020 374052 287026
rect 374000 286962 374052 286968
rect 374656 284306 374684 307838
rect 389376 305946 389404 307906
rect 399024 307828 399076 307834
rect 399024 307770 399076 307776
rect 399036 305946 399064 307770
rect 389376 305918 389712 305946
rect 399036 305918 399372 305946
rect 379624 305238 380052 305266
rect 378046 296304 378102 296313
rect 378046 296239 378102 296248
rect 378060 286890 378088 296239
rect 378048 286884 378100 286890
rect 378048 286826 378100 286832
rect 374644 284300 374696 284306
rect 374644 284242 374696 284248
rect 379624 284170 379652 305238
rect 399496 286770 399524 307906
rect 400864 307828 400916 307834
rect 400864 307770 400916 307776
rect 399372 286742 399524 286770
rect 379716 286062 380052 286090
rect 389712 286062 390048 286090
rect 379716 284306 379744 286062
rect 379704 284300 379756 284306
rect 379704 284242 379756 284248
rect 352012 284164 352064 284170
rect 352012 284106 352064 284112
rect 361672 284164 361724 284170
rect 361672 284106 361724 284112
rect 373264 284164 373316 284170
rect 373264 284106 373316 284112
rect 379612 284164 379664 284170
rect 379612 284106 379664 284112
rect 390020 284102 390048 286062
rect 400876 284102 400904 307770
rect 408052 305932 408080 307974
rect 417700 307964 417752 307970
rect 417700 307906 417752 307912
rect 417712 305932 417740 307906
rect 428556 307896 428608 307902
rect 428556 307838 428608 307844
rect 427360 307828 427412 307834
rect 427360 307770 427412 307776
rect 428464 307828 428516 307834
rect 428464 307770 428516 307776
rect 427372 305932 427400 307770
rect 405646 296304 405702 296313
rect 405646 296239 405702 296248
rect 401598 295624 401654 295633
rect 401598 295559 401654 295568
rect 401612 286958 401640 295559
rect 405660 287026 405688 296239
rect 405648 287020 405700 287026
rect 405648 286962 405700 286968
rect 401600 286952 401652 286958
rect 401600 286894 401652 286900
rect 427728 286816 427780 286822
rect 427386 286764 427728 286770
rect 427386 286758 427780 286764
rect 427386 286742 427768 286758
rect 408052 284170 408080 286076
rect 417712 284170 417740 286076
rect 428476 284170 428504 307770
rect 428568 286822 428596 307838
rect 428660 287706 428688 307974
rect 456064 307964 456116 307970
rect 456064 307906 456116 307912
rect 473544 307964 473596 307970
rect 473544 307906 473596 307912
rect 483480 307964 483532 307970
rect 483480 307906 483532 307912
rect 445668 307896 445720 307902
rect 445668 307838 445720 307844
rect 445680 305932 445708 307838
rect 455328 307828 455380 307834
rect 455328 307770 455380 307776
rect 455340 305932 455368 307770
rect 434824 305238 436034 305266
rect 434626 296304 434682 296313
rect 434626 296239 434682 296248
rect 429198 295624 429254 295633
rect 429198 295559 429254 295568
rect 428648 287700 428700 287706
rect 428648 287642 428700 287648
rect 429212 286890 429240 295559
rect 434640 286958 434668 296239
rect 434628 286952 434680 286958
rect 434628 286894 434680 286900
rect 429200 286884 429252 286890
rect 429200 286826 429252 286832
rect 428556 286816 428608 286822
rect 428556 286758 428608 286764
rect 434824 284170 434852 305238
rect 435732 287700 435784 287706
rect 435732 287642 435784 287648
rect 435744 286770 435772 287642
rect 456076 287054 456104 307906
rect 464344 307896 464396 307902
rect 464344 307838 464396 307844
rect 456156 307828 456208 307834
rect 456156 307770 456208 307776
rect 455800 287026 456104 287054
rect 455800 286770 455828 287026
rect 435744 286742 436034 286770
rect 455354 286742 455828 286770
rect 408040 284164 408092 284170
rect 408040 284106 408092 284112
rect 417700 284164 417752 284170
rect 417700 284106 417752 284112
rect 428464 284164 428516 284170
rect 428464 284106 428516 284112
rect 434812 284164 434864 284170
rect 434812 284106 434864 284112
rect 445680 284102 445708 286076
rect 456168 284102 456196 307770
rect 464356 305946 464384 307838
rect 464048 305918 464384 305946
rect 473556 305946 473584 307906
rect 483204 307828 483256 307834
rect 483204 307770 483256 307776
rect 483216 305946 483244 307770
rect 473556 305918 473708 305946
rect 483216 305918 483368 305946
rect 462226 296304 462282 296313
rect 462226 296239 462282 296248
rect 458178 295624 458234 295633
rect 458178 295559 458234 295568
rect 458192 287026 458220 295559
rect 458180 287020 458232 287026
rect 458180 286962 458232 286968
rect 462240 286890 462268 296239
rect 462228 286884 462280 286890
rect 462228 286826 462280 286832
rect 483492 286770 483520 307906
rect 483664 307896 483716 307902
rect 483664 307838 483716 307844
rect 483676 287434 483704 307838
rect 485044 307828 485096 307834
rect 485044 307770 485096 307776
rect 483664 287428 483716 287434
rect 483664 287370 483716 287376
rect 483368 286742 483520 286770
rect 463712 286062 464048 286090
rect 473708 286062 474044 286090
rect 463712 284170 463740 286062
rect 474016 284170 474044 286062
rect 485056 284170 485084 307770
rect 489826 296304 489882 296313
rect 489826 296239 489882 296248
rect 485778 295624 485834 295633
rect 485778 295559 485834 295568
rect 485792 286958 485820 295559
rect 489840 287026 489868 296239
rect 489828 287020 489880 287026
rect 489828 286962 489880 286968
rect 485780 286952 485832 286958
rect 485780 286894 485832 286900
rect 463700 284164 463752 284170
rect 463700 284106 463752 284112
rect 474004 284164 474056 284170
rect 474004 284106 474056 284112
rect 485044 284164 485096 284170
rect 485044 284106 485096 284112
rect 333704 284096 333756 284102
rect 333704 284038 333756 284044
rect 344284 284096 344336 284102
rect 344284 284038 344336 284044
rect 390008 284096 390060 284102
rect 390008 284038 390060 284044
rect 400864 284096 400916 284102
rect 400864 284038 400916 284044
rect 445668 284096 445720 284102
rect 445668 284038 445720 284044
rect 456156 284096 456208 284102
rect 456156 284038 456208 284044
rect 296352 280424 296404 280430
rect 296352 280366 296404 280372
rect 316776 280424 316828 280430
rect 316776 280366 316828 280372
rect 408040 280424 408092 280430
rect 408040 280366 408092 280372
rect 428648 280424 428700 280430
rect 428648 280366 428700 280372
rect 277676 280356 277728 280362
rect 277676 280298 277728 280304
rect 287520 280356 287572 280362
rect 287520 280298 287572 280304
rect 268016 280288 268068 280294
rect 268016 280230 268068 280236
rect 268028 278868 268056 280230
rect 277688 278868 277716 280298
rect 287336 280220 287388 280226
rect 287336 280162 287388 280168
rect 287348 278868 287376 280162
rect 262220 277432 262272 277438
rect 262220 277374 262272 277380
rect 266268 277432 266320 277438
rect 266268 277374 266320 277380
rect 262232 268569 262260 277374
rect 266280 269249 266308 277374
rect 266266 269240 266322 269249
rect 266266 269175 266322 269184
rect 262218 268560 262274 268569
rect 262218 268495 262274 268504
rect 287532 259706 287560 280298
rect 287704 280288 287756 280294
rect 287704 280230 287756 280236
rect 287716 261322 287744 280230
rect 289084 280220 289136 280226
rect 289084 280162 289136 280168
rect 287704 261316 287756 261322
rect 287704 261258 287756 261264
rect 287362 259678 287560 259706
rect 249708 256624 249760 256630
rect 249708 256566 249760 256572
rect 260196 256624 260248 256630
rect 260196 256566 260248 256572
rect 261484 256624 261536 256630
rect 261484 256566 261536 256572
rect 268028 256562 268056 259148
rect 277688 256562 277716 259148
rect 289096 256562 289124 280162
rect 296364 278882 296392 280366
rect 305368 280356 305420 280362
rect 305368 280298 305420 280304
rect 296056 278854 296392 278882
rect 305380 278882 305408 280298
rect 315488 280288 315540 280294
rect 315488 280230 315540 280236
rect 315028 280220 315080 280226
rect 315028 280162 315080 280168
rect 315040 278882 315068 280162
rect 305380 278854 305716 278882
rect 315040 278854 315376 278882
rect 289820 277500 289872 277506
rect 289820 277442 289872 277448
rect 293868 277500 293920 277506
rect 293868 277442 293920 277448
rect 289832 268569 289860 277442
rect 293880 269249 293908 277442
rect 293866 269240 293922 269249
rect 293866 269175 293922 269184
rect 289818 268560 289874 268569
rect 289818 268495 289874 268504
rect 295708 261316 295760 261322
rect 295708 261258 295760 261264
rect 295720 259706 295748 261258
rect 315500 259706 315528 280230
rect 316684 280220 316736 280226
rect 316684 280162 316736 280168
rect 295720 259678 296056 259706
rect 315376 259678 315528 259706
rect 305716 259134 306052 259162
rect 306024 256562 306052 259134
rect 316696 256562 316724 280162
rect 316788 261458 316816 280366
rect 345664 280356 345716 280362
rect 345664 280298 345716 280304
rect 361672 280356 361724 280362
rect 361672 280298 361724 280304
rect 371516 280356 371568 280362
rect 371516 280298 371568 280304
rect 389364 280356 389416 280362
rect 389364 280298 389416 280304
rect 399484 280356 399536 280362
rect 399484 280298 399536 280304
rect 333704 280288 333756 280294
rect 333704 280230 333756 280236
rect 333716 278868 333744 280230
rect 343364 280220 343416 280226
rect 343364 280162 343416 280168
rect 344284 280220 344336 280226
rect 344284 280162 344336 280168
rect 343376 278868 343404 280162
rect 323044 278310 324070 278338
rect 317420 277432 317472 277438
rect 317420 277374 317472 277380
rect 322848 277432 322900 277438
rect 322848 277374 322900 277380
rect 317432 268569 317460 277374
rect 322860 269249 322888 277374
rect 322846 269240 322902 269249
rect 322846 269175 322902 269184
rect 317418 268560 317474 268569
rect 317418 268495 317474 268504
rect 316776 261452 316828 261458
rect 316776 261394 316828 261400
rect 323044 256562 323072 278310
rect 323676 261452 323728 261458
rect 323676 261394 323728 261400
rect 323688 259706 323716 261394
rect 323688 259678 324070 259706
rect 343390 259418 343680 259434
rect 343390 259412 343692 259418
rect 343390 259406 343640 259412
rect 343640 259354 343692 259360
rect 238852 256556 238904 256562
rect 238852 256498 238904 256504
rect 268016 256556 268068 256562
rect 268016 256498 268068 256504
rect 277676 256556 277728 256562
rect 277676 256498 277728 256504
rect 289084 256556 289136 256562
rect 289084 256498 289136 256504
rect 306012 256556 306064 256562
rect 306012 256498 306064 256504
rect 316684 256556 316736 256562
rect 316684 256498 316736 256504
rect 323032 256556 323084 256562
rect 323032 256498 323084 256504
rect 333716 256494 333744 259148
rect 344296 256494 344324 280162
rect 345020 277500 345072 277506
rect 345020 277442 345072 277448
rect 345032 268569 345060 277442
rect 345018 268560 345074 268569
rect 345018 268495 345074 268504
rect 345676 259418 345704 280298
rect 352012 280288 352064 280294
rect 352012 280230 352064 280236
rect 352024 278868 352052 280230
rect 361684 278868 361712 280298
rect 371332 280220 371384 280226
rect 371332 280162 371384 280168
rect 371344 278868 371372 280162
rect 350448 277500 350500 277506
rect 350448 277442 350500 277448
rect 350460 269249 350488 277442
rect 350446 269240 350502 269249
rect 350446 269175 350502 269184
rect 371528 259706 371556 280298
rect 374644 280288 374696 280294
rect 374644 280230 374696 280236
rect 373264 280220 373316 280226
rect 373264 280162 373316 280168
rect 371358 259678 371556 259706
rect 345664 259412 345716 259418
rect 345664 259354 345716 259360
rect 352024 256562 352052 259148
rect 361684 256562 361712 259148
rect 373276 256562 373304 280162
rect 374000 277432 374052 277438
rect 374000 277374 374052 277380
rect 374012 269113 374040 277374
rect 373998 269104 374054 269113
rect 373998 269039 374054 269048
rect 374656 256698 374684 280230
rect 389376 278882 389404 280298
rect 399024 280220 399076 280226
rect 399024 280162 399076 280168
rect 399036 278882 399064 280162
rect 389376 278854 389712 278882
rect 399036 278854 399372 278882
rect 379624 278310 380052 278338
rect 378048 277568 378100 277574
rect 378048 277510 378100 277516
rect 378060 269249 378088 277510
rect 378046 269240 378102 269249
rect 378046 269175 378102 269184
rect 374644 256692 374696 256698
rect 374644 256634 374696 256640
rect 379624 256562 379652 278310
rect 399496 259706 399524 280298
rect 400864 280220 400916 280226
rect 400864 280162 400916 280168
rect 399372 259678 399524 259706
rect 379716 259134 380052 259162
rect 389712 259134 390048 259162
rect 379716 256698 379744 259134
rect 379704 256692 379756 256698
rect 379704 256634 379756 256640
rect 352012 256556 352064 256562
rect 352012 256498 352064 256504
rect 361672 256556 361724 256562
rect 361672 256498 361724 256504
rect 373264 256556 373316 256562
rect 373264 256498 373316 256504
rect 379612 256556 379664 256562
rect 379612 256498 379664 256504
rect 390020 256494 390048 259134
rect 400876 256494 400904 280162
rect 408052 278868 408080 280366
rect 417700 280356 417752 280362
rect 417700 280298 417752 280304
rect 417712 278868 417740 280298
rect 428464 280288 428516 280294
rect 428464 280230 428516 280236
rect 427360 280220 427412 280226
rect 427360 280162 427412 280168
rect 427372 278868 427400 280162
rect 401600 277500 401652 277506
rect 401600 277442 401652 277448
rect 401612 268569 401640 277442
rect 405648 277432 405700 277438
rect 405648 277374 405700 277380
rect 405660 269249 405688 277374
rect 405646 269240 405702 269249
rect 405646 269175 405702 269184
rect 401598 268560 401654 268569
rect 401598 268495 401654 268504
rect 428476 267734 428504 280230
rect 428556 280220 428608 280226
rect 428556 280162 428608 280168
rect 427832 267706 428504 267734
rect 427832 259434 427860 267706
rect 427386 259406 427860 259434
rect 408052 256562 408080 259148
rect 417712 256562 417740 259148
rect 428568 256562 428596 280162
rect 428660 261526 428688 280366
rect 456156 280356 456208 280362
rect 456156 280298 456208 280304
rect 473360 280356 473412 280362
rect 473360 280298 473412 280304
rect 483480 280356 483532 280362
rect 483480 280298 483532 280304
rect 445668 280288 445720 280294
rect 445668 280230 445720 280236
rect 445680 278868 445708 280230
rect 455328 280220 455380 280226
rect 455328 280162 455380 280168
rect 456064 280220 456116 280226
rect 456064 280162 456116 280168
rect 455340 278868 455368 280162
rect 434824 278310 436034 278338
rect 429200 277568 429252 277574
rect 429200 277510 429252 277516
rect 429212 268569 429240 277510
rect 434628 277500 434680 277506
rect 434628 277442 434680 277448
rect 434640 269249 434668 277442
rect 434626 269240 434682 269249
rect 434626 269175 434682 269184
rect 429198 268560 429254 268569
rect 429198 268495 429254 268504
rect 428648 261520 428700 261526
rect 428648 261462 428700 261468
rect 434824 256562 434852 278310
rect 455696 263492 455748 263498
rect 455696 263434 455748 263440
rect 435732 261520 435784 261526
rect 435732 261462 435784 261468
rect 435744 259706 435772 261462
rect 455708 259706 455736 263434
rect 435744 259678 436034 259706
rect 455354 259678 455736 259706
rect 408040 256556 408092 256562
rect 408040 256498 408092 256504
rect 417700 256556 417752 256562
rect 417700 256498 417752 256504
rect 428556 256556 428608 256562
rect 428556 256498 428608 256504
rect 434812 256556 434864 256562
rect 434812 256498 434864 256504
rect 445680 256494 445708 259148
rect 456076 256494 456104 280162
rect 456168 263498 456196 280298
rect 464344 280288 464396 280294
rect 464344 280230 464396 280236
rect 464356 278882 464384 280230
rect 464048 278854 464384 278882
rect 473372 278882 473400 280298
rect 483020 280220 483072 280226
rect 483020 280162 483072 280168
rect 483032 278882 483060 280162
rect 473372 278854 473708 278882
rect 483032 278854 483368 278882
rect 462228 277568 462280 277574
rect 462228 277510 462280 277516
rect 458180 277432 458232 277438
rect 458180 277374 458232 277380
rect 458192 268569 458220 277374
rect 462240 269249 462268 277510
rect 462226 269240 462282 269249
rect 462226 269175 462282 269184
rect 458178 268560 458234 268569
rect 458178 268495 458234 268504
rect 456156 263492 456208 263498
rect 456156 263434 456208 263440
rect 483492 259706 483520 280298
rect 483664 280288 483716 280294
rect 483664 280230 483716 280236
rect 483676 262206 483704 280230
rect 485044 280220 485096 280226
rect 485044 280162 485096 280168
rect 483664 262200 483716 262206
rect 483664 262142 483716 262148
rect 483368 259678 483520 259706
rect 463804 259134 464048 259162
rect 473708 259134 474044 259162
rect 463804 256562 463832 259134
rect 474016 256562 474044 259134
rect 485056 256562 485084 280162
rect 485780 277500 485832 277506
rect 485780 277442 485832 277448
rect 485792 268569 485820 277442
rect 489828 277432 489880 277438
rect 489828 277374 489880 277380
rect 489840 269249 489868 277374
rect 489826 269240 489882 269249
rect 489826 269175 489882 269184
rect 485778 268560 485834 268569
rect 485778 268495 485834 268504
rect 463792 256556 463844 256562
rect 463792 256498 463844 256504
rect 474004 256556 474056 256562
rect 474004 256498 474056 256504
rect 485044 256556 485096 256562
rect 485044 256498 485096 256504
rect 333704 256488 333756 256494
rect 333704 256430 333756 256436
rect 344284 256488 344336 256494
rect 344284 256430 344336 256436
rect 390008 256488 390060 256494
rect 390008 256430 390060 256436
rect 400864 256488 400916 256494
rect 400864 256430 400916 256436
rect 445668 256488 445720 256494
rect 445668 256430 445720 256436
rect 456064 256488 456116 256494
rect 456064 256430 456116 256436
rect 296352 254176 296404 254182
rect 296352 254118 296404 254124
rect 316776 254176 316828 254182
rect 316776 254118 316828 254124
rect 260196 254108 260248 254114
rect 260196 254050 260248 254056
rect 277676 254108 277728 254114
rect 277676 254050 277728 254056
rect 287520 254108 287572 254114
rect 287520 254050 287572 254056
rect 249708 254040 249760 254046
rect 249708 253982 249760 253988
rect 249720 251940 249748 253982
rect 259368 253972 259420 253978
rect 259368 253914 259420 253920
rect 260104 253972 260156 253978
rect 260104 253914 260156 253920
rect 259380 251940 259408 253914
rect 238668 251252 238720 251258
rect 238668 251194 238720 251200
rect 238864 251246 240074 251274
rect 238680 242321 238708 251194
rect 238666 242312 238722 242321
rect 238666 242247 238722 242256
rect 238864 230314 238892 251246
rect 259736 235408 259788 235414
rect 259736 235350 259788 235356
rect 239772 233572 239824 233578
rect 239772 233514 239824 233520
rect 239784 232778 239812 233514
rect 259748 232778 259776 235350
rect 239784 232750 240074 232778
rect 259394 232750 259776 232778
rect 238852 230308 238904 230314
rect 238852 230250 238904 230256
rect 249720 230246 249748 232084
rect 260116 230246 260144 253914
rect 260208 235414 260236 254050
rect 268016 254040 268068 254046
rect 268016 253982 268068 253988
rect 268028 251940 268056 253982
rect 277688 251940 277716 254050
rect 287336 253972 287388 253978
rect 287336 253914 287388 253920
rect 287348 251940 287376 253914
rect 266266 242312 266322 242321
rect 266266 242247 266322 242256
rect 262218 241632 262274 241641
rect 262218 241567 262274 241576
rect 260196 235408 260248 235414
rect 260196 235350 260248 235356
rect 262232 233238 262260 241567
rect 266280 233238 266308 242247
rect 262220 233232 262272 233238
rect 262220 233174 262272 233180
rect 266268 233232 266320 233238
rect 266268 233174 266320 233180
rect 287532 232778 287560 254050
rect 287704 254040 287756 254046
rect 287704 253982 287756 253988
rect 287716 233578 287744 253982
rect 289084 253972 289136 253978
rect 289084 253914 289136 253920
rect 287704 233572 287756 233578
rect 287704 233514 287756 233520
rect 287362 232750 287560 232778
rect 268028 230314 268056 232084
rect 277688 230314 277716 232084
rect 289096 230314 289124 253914
rect 296364 251954 296392 254118
rect 305368 254108 305420 254114
rect 305368 254050 305420 254056
rect 296056 251926 296392 251954
rect 305380 251954 305408 254050
rect 315488 254040 315540 254046
rect 315488 253982 315540 253988
rect 315028 253972 315080 253978
rect 315028 253914 315080 253920
rect 315040 251954 315068 253914
rect 305380 251926 305716 251954
rect 315040 251926 315376 251954
rect 289820 251252 289872 251258
rect 289820 251194 289872 251200
rect 293868 251252 293920 251258
rect 293868 251194 293920 251200
rect 289832 241641 289860 251194
rect 293880 242321 293908 251194
rect 293866 242312 293922 242321
rect 293866 242247 293922 242256
rect 289818 241632 289874 241641
rect 289818 241567 289874 241576
rect 295708 233572 295760 233578
rect 295708 233514 295760 233520
rect 295720 232778 295748 233514
rect 315500 232778 315528 253982
rect 316684 253972 316736 253978
rect 316684 253914 316736 253920
rect 295720 232750 296056 232778
rect 315376 232750 315528 232778
rect 305716 232070 306052 232098
rect 306024 230314 306052 232070
rect 316696 230314 316724 253914
rect 316788 233442 316816 254118
rect 345664 254108 345716 254114
rect 345664 254050 345716 254056
rect 361672 254108 361724 254114
rect 361672 254050 361724 254056
rect 371516 254108 371568 254114
rect 371516 254050 371568 254056
rect 389364 254108 389416 254114
rect 389364 254050 389416 254056
rect 399484 254108 399536 254114
rect 399484 254050 399536 254056
rect 417700 254108 417752 254114
rect 417700 254050 417752 254056
rect 428556 254108 428608 254114
rect 428556 254050 428608 254056
rect 445668 254108 445720 254114
rect 445668 254050 445720 254056
rect 456064 254108 456116 254114
rect 456064 254050 456116 254056
rect 473360 254108 473412 254114
rect 473360 254050 473412 254056
rect 483480 254108 483532 254114
rect 483480 254050 483532 254056
rect 333704 254040 333756 254046
rect 333704 253982 333756 253988
rect 333716 251940 333744 253982
rect 343364 253972 343416 253978
rect 343364 253914 343416 253920
rect 344284 253972 344336 253978
rect 344284 253914 344336 253920
rect 343376 251940 343404 253914
rect 323044 251246 324070 251274
rect 322846 242312 322902 242321
rect 322846 242247 322902 242256
rect 317418 241632 317474 241641
rect 317418 241567 317474 241576
rect 316776 233436 316828 233442
rect 316776 233378 316828 233384
rect 317432 233238 317460 241567
rect 322860 233238 322888 242247
rect 317420 233232 317472 233238
rect 317420 233174 317472 233180
rect 322848 233232 322900 233238
rect 322848 233174 322900 233180
rect 323044 230314 323072 251246
rect 323676 233436 323728 233442
rect 323676 233378 323728 233384
rect 323688 232778 323716 233378
rect 323688 232750 324070 232778
rect 343390 232762 343680 232778
rect 343390 232756 343692 232762
rect 343390 232750 343640 232756
rect 343640 232698 343692 232704
rect 268016 230308 268068 230314
rect 268016 230250 268068 230256
rect 277676 230308 277728 230314
rect 277676 230250 277728 230256
rect 289084 230308 289136 230314
rect 289084 230250 289136 230256
rect 306012 230308 306064 230314
rect 306012 230250 306064 230256
rect 316684 230308 316736 230314
rect 316684 230250 316736 230256
rect 323032 230308 323084 230314
rect 323032 230250 323084 230256
rect 333716 230246 333744 232084
rect 344296 230246 344324 253914
rect 345020 251252 345072 251258
rect 345020 251194 345072 251200
rect 345032 241641 345060 251194
rect 345018 241632 345074 241641
rect 345018 241567 345074 241576
rect 345676 232762 345704 254050
rect 352012 254040 352064 254046
rect 352012 253982 352064 253988
rect 352024 251940 352052 253982
rect 361684 251940 361712 254050
rect 371332 253972 371384 253978
rect 371332 253914 371384 253920
rect 371344 251940 371372 253914
rect 350448 251252 350500 251258
rect 350448 251194 350500 251200
rect 350460 242321 350488 251194
rect 350446 242312 350502 242321
rect 350446 242247 350502 242256
rect 371528 232778 371556 254050
rect 374644 254040 374696 254046
rect 374644 253982 374696 253988
rect 373264 253972 373316 253978
rect 373264 253914 373316 253920
rect 345664 232756 345716 232762
rect 371358 232750 371556 232778
rect 345664 232698 345716 232704
rect 352024 230314 352052 232084
rect 361684 230314 361712 232084
rect 373276 230314 373304 253914
rect 373998 241632 374054 241641
rect 373998 241567 374054 241576
rect 374012 233238 374040 241567
rect 374000 233232 374052 233238
rect 374000 233174 374052 233180
rect 374656 230450 374684 253982
rect 389376 251954 389404 254050
rect 399024 253972 399076 253978
rect 399024 253914 399076 253920
rect 399036 251954 399064 253914
rect 389376 251926 389712 251954
rect 399036 251926 399372 251954
rect 378048 251320 378100 251326
rect 378048 251262 378100 251268
rect 378060 242321 378088 251262
rect 379624 251246 380052 251274
rect 378046 242312 378102 242321
rect 378046 242247 378102 242256
rect 374644 230444 374696 230450
rect 374644 230386 374696 230392
rect 379624 230314 379652 251246
rect 399496 232778 399524 254050
rect 408040 254040 408092 254046
rect 408040 253982 408092 253988
rect 400864 253972 400916 253978
rect 400864 253914 400916 253920
rect 399372 232750 399524 232778
rect 379716 232070 380052 232098
rect 389712 232070 390048 232098
rect 379716 230450 379744 232070
rect 379704 230444 379756 230450
rect 379704 230386 379756 230392
rect 352012 230308 352064 230314
rect 352012 230250 352064 230256
rect 361672 230308 361724 230314
rect 361672 230250 361724 230256
rect 373264 230308 373316 230314
rect 373264 230250 373316 230256
rect 379612 230308 379664 230314
rect 379612 230250 379664 230256
rect 390020 230246 390048 232070
rect 400876 230246 400904 253914
rect 408052 251940 408080 253982
rect 417712 251940 417740 254050
rect 427360 253972 427412 253978
rect 427360 253914 427412 253920
rect 428464 253972 428516 253978
rect 428464 253914 428516 253920
rect 427372 251940 427400 253914
rect 401600 251252 401652 251258
rect 401600 251194 401652 251200
rect 401612 241641 401640 251194
rect 405646 242312 405702 242321
rect 405646 242247 405702 242256
rect 401598 241632 401654 241641
rect 401598 241567 401654 241576
rect 405660 233238 405688 242247
rect 405648 233232 405700 233238
rect 405648 233174 405700 233180
rect 427728 233164 427780 233170
rect 427728 233106 427780 233112
rect 427740 232778 427768 233106
rect 427386 232750 427768 232778
rect 408052 230314 408080 232084
rect 417712 230314 417740 232084
rect 428476 230314 428504 253914
rect 428568 233170 428596 254050
rect 428648 254040 428700 254046
rect 428648 253982 428700 253988
rect 428660 233918 428688 253982
rect 445680 251940 445708 254050
rect 455328 253972 455380 253978
rect 455328 253914 455380 253920
rect 455340 251940 455368 253914
rect 429200 251320 429252 251326
rect 429200 251262 429252 251268
rect 429212 241641 429240 251262
rect 434628 251252 434680 251258
rect 434628 251194 434680 251200
rect 434824 251246 436034 251274
rect 434640 242321 434668 251194
rect 434626 242312 434682 242321
rect 434626 242247 434682 242256
rect 429198 241632 429254 241641
rect 429198 241567 429254 241576
rect 428648 233912 428700 233918
rect 428648 233854 428700 233860
rect 428556 233164 428608 233170
rect 428556 233106 428608 233112
rect 434824 230314 434852 251246
rect 456076 238754 456104 254050
rect 464344 254040 464396 254046
rect 464344 253982 464396 253988
rect 456156 253972 456208 253978
rect 456156 253914 456208 253920
rect 455800 238726 456104 238754
rect 435732 233912 435784 233918
rect 435732 233854 435784 233860
rect 435744 232778 435772 233854
rect 455800 232778 455828 238726
rect 435744 232750 436034 232778
rect 455354 232750 455828 232778
rect 408040 230308 408092 230314
rect 408040 230250 408092 230256
rect 417700 230308 417752 230314
rect 417700 230250 417752 230256
rect 428464 230308 428516 230314
rect 428464 230250 428516 230256
rect 434812 230308 434864 230314
rect 434812 230250 434864 230256
rect 445680 230246 445708 232084
rect 456168 230246 456196 253914
rect 464356 251954 464384 253982
rect 464048 251926 464384 251954
rect 473372 251954 473400 254050
rect 483020 253972 483072 253978
rect 483020 253914 483072 253920
rect 483032 251954 483060 253914
rect 473372 251926 473708 251954
rect 483032 251926 483368 251954
rect 462226 242312 462282 242321
rect 462226 242247 462282 242256
rect 458178 241632 458234 241641
rect 458178 241567 458234 241576
rect 458192 233238 458220 241567
rect 462240 233238 462268 242247
rect 458180 233232 458232 233238
rect 458180 233174 458232 233180
rect 462228 233232 462280 233238
rect 462228 233174 462280 233180
rect 483492 232778 483520 254050
rect 483664 254040 483716 254046
rect 483664 253982 483716 253988
rect 483676 233442 483704 253982
rect 485044 253972 485096 253978
rect 485044 253914 485096 253920
rect 483664 233436 483716 233442
rect 483664 233378 483716 233384
rect 483368 232750 483520 232778
rect 463712 232070 464048 232098
rect 473708 232070 474044 232098
rect 463712 230314 463740 232070
rect 474016 230314 474044 232070
rect 485056 230314 485084 253914
rect 485780 251252 485832 251258
rect 485780 251194 485832 251200
rect 489828 251252 489880 251258
rect 489828 251194 489880 251200
rect 485792 241641 485820 251194
rect 489840 242321 489868 251194
rect 489826 242312 489882 242321
rect 489826 242247 489882 242256
rect 485778 241632 485834 241641
rect 485778 241567 485834 241576
rect 463700 230308 463752 230314
rect 463700 230250 463752 230256
rect 474004 230308 474056 230314
rect 474004 230250 474056 230256
rect 485044 230308 485096 230314
rect 485044 230250 485096 230256
rect 249708 230240 249760 230246
rect 249708 230182 249760 230188
rect 260104 230240 260156 230246
rect 260104 230182 260156 230188
rect 333704 230240 333756 230246
rect 333704 230182 333756 230188
rect 344284 230240 344336 230246
rect 344284 230182 344336 230188
rect 390008 230240 390060 230246
rect 390008 230182 390060 230188
rect 400864 230240 400916 230246
rect 400864 230182 400916 230188
rect 445668 230240 445720 230246
rect 445668 230182 445720 230188
rect 456156 230240 456208 230246
rect 456156 230182 456208 230188
rect 261484 226636 261536 226642
rect 261484 226578 261536 226584
rect 249708 226500 249760 226506
rect 249708 226442 249760 226448
rect 260196 226500 260248 226506
rect 260196 226442 260248 226448
rect 249720 224876 249748 226442
rect 259368 226432 259420 226438
rect 259368 226374 259420 226380
rect 259380 224876 259408 226374
rect 260104 226364 260156 226370
rect 260104 226306 260156 226312
rect 238864 224318 240074 224346
rect 238666 215248 238722 215257
rect 238666 215183 238722 215192
rect 238680 205562 238708 215183
rect 238668 205556 238720 205562
rect 238668 205498 238720 205504
rect 238864 202706 238892 224318
rect 239772 207800 239824 207806
rect 239772 207742 239824 207748
rect 239784 205714 239812 207742
rect 259736 207392 259788 207398
rect 259736 207334 259788 207340
rect 259748 205714 259776 207334
rect 239784 205686 240074 205714
rect 259394 205686 259776 205714
rect 249536 205142 249734 205170
rect 238852 202700 238904 202706
rect 238852 202642 238904 202648
rect 249536 202638 249564 205142
rect 260116 202638 260144 226306
rect 260208 207398 260236 226442
rect 260196 207392 260248 207398
rect 260196 207334 260248 207340
rect 249524 202632 249576 202638
rect 249524 202574 249576 202580
rect 260104 202632 260156 202638
rect 260104 202574 260156 202580
rect 260196 200320 260248 200326
rect 260196 200262 260248 200268
rect 249708 200252 249760 200258
rect 249708 200194 249760 200200
rect 249720 197948 249748 200194
rect 259368 200184 259420 200190
rect 259368 200126 259420 200132
rect 260104 200184 260156 200190
rect 260104 200126 260156 200132
rect 259380 197948 259408 200126
rect 238864 197254 240074 197282
rect 238666 188320 238722 188329
rect 238666 188255 238722 188264
rect 238680 179314 238708 188255
rect 238668 179308 238720 179314
rect 238668 179250 238720 179256
rect 238864 176526 238892 197254
rect 259736 185632 259788 185638
rect 259736 185574 259788 185580
rect 239772 179920 239824 179926
rect 239772 179862 239824 179868
rect 239784 178786 239812 179862
rect 259748 178786 259776 185574
rect 239784 178758 240074 178786
rect 259394 178758 259776 178786
rect 249720 176594 249748 178092
rect 260116 176594 260144 200126
rect 260208 185638 260236 200262
rect 260196 185632 260248 185638
rect 260196 185574 260248 185580
rect 261496 176594 261524 226578
rect 296352 226568 296404 226574
rect 296352 226510 296404 226516
rect 316776 226568 316828 226574
rect 316776 226510 316828 226516
rect 408040 226568 408092 226574
rect 408040 226510 408092 226516
rect 428648 226568 428700 226574
rect 428648 226510 428700 226516
rect 277676 226500 277728 226506
rect 277676 226442 277728 226448
rect 287520 226500 287572 226506
rect 287520 226442 287572 226448
rect 268016 226432 268068 226438
rect 268016 226374 268068 226380
rect 268028 224876 268056 226374
rect 277688 224876 277716 226442
rect 287336 226364 287388 226370
rect 287336 226306 287388 226312
rect 287348 224876 287376 226306
rect 266266 215248 266322 215257
rect 266266 215183 266322 215192
rect 262218 214568 262274 214577
rect 262218 214503 262274 214512
rect 262232 205630 262260 214503
rect 266280 205630 266308 215183
rect 287532 205714 287560 226442
rect 287704 226432 287756 226438
rect 287704 226374 287756 226380
rect 287716 207194 287744 226374
rect 289084 226364 289136 226370
rect 289084 226306 289136 226312
rect 287704 207188 287756 207194
rect 287704 207130 287756 207136
rect 287362 205686 287560 205714
rect 262220 205624 262272 205630
rect 262220 205566 262272 205572
rect 266268 205624 266320 205630
rect 266268 205566 266320 205572
rect 268028 202706 268056 205020
rect 277688 202706 277716 205020
rect 289096 202706 289124 226306
rect 296364 224890 296392 226510
rect 305368 226500 305420 226506
rect 305368 226442 305420 226448
rect 296056 224862 296392 224890
rect 305380 224890 305408 226442
rect 315488 226432 315540 226438
rect 315488 226374 315540 226380
rect 315028 226364 315080 226370
rect 315028 226306 315080 226312
rect 315040 224890 315068 226306
rect 305380 224862 305716 224890
rect 315040 224862 315376 224890
rect 293866 215248 293922 215257
rect 293866 215183 293922 215192
rect 289818 214568 289874 214577
rect 289818 214503 289874 214512
rect 289832 205562 289860 214503
rect 293880 205562 293908 215183
rect 295708 207188 295760 207194
rect 295708 207130 295760 207136
rect 295720 205714 295748 207130
rect 315500 205714 315528 226374
rect 316684 226364 316736 226370
rect 316684 226306 316736 226312
rect 295720 205686 296056 205714
rect 315376 205686 315528 205714
rect 289820 205556 289872 205562
rect 289820 205498 289872 205504
rect 293868 205556 293920 205562
rect 293868 205498 293920 205504
rect 305716 205006 306052 205034
rect 306024 202706 306052 205006
rect 316696 202706 316724 226306
rect 316788 207398 316816 226510
rect 345664 226500 345716 226506
rect 345664 226442 345716 226448
rect 361672 226500 361724 226506
rect 361672 226442 361724 226448
rect 371516 226500 371568 226506
rect 371516 226442 371568 226448
rect 389364 226500 389416 226506
rect 389364 226442 389416 226448
rect 399484 226500 399536 226506
rect 399484 226442 399536 226448
rect 333704 226432 333756 226438
rect 333704 226374 333756 226380
rect 333716 224876 333744 226374
rect 343364 226364 343416 226370
rect 343364 226306 343416 226312
rect 344284 226364 344336 226370
rect 344284 226306 344336 226312
rect 343376 224876 343404 226306
rect 323044 224318 324070 224346
rect 322846 215248 322902 215257
rect 322846 215183 322902 215192
rect 317418 214568 317474 214577
rect 317418 214503 317474 214512
rect 316776 207392 316828 207398
rect 316776 207334 316828 207340
rect 317432 205630 317460 214503
rect 322860 205630 322888 215183
rect 317420 205624 317472 205630
rect 317420 205566 317472 205572
rect 322848 205624 322900 205630
rect 322848 205566 322900 205572
rect 323044 202706 323072 224318
rect 323676 207392 323728 207398
rect 323676 207334 323728 207340
rect 323688 205714 323716 207334
rect 323688 205686 324070 205714
rect 343640 205488 343692 205494
rect 343390 205436 343640 205442
rect 343390 205430 343692 205436
rect 343390 205414 343680 205430
rect 333730 205006 333928 205034
rect 268016 202700 268068 202706
rect 268016 202642 268068 202648
rect 277676 202700 277728 202706
rect 277676 202642 277728 202648
rect 289084 202700 289136 202706
rect 289084 202642 289136 202648
rect 306012 202700 306064 202706
rect 306012 202642 306064 202648
rect 316684 202700 316736 202706
rect 316684 202642 316736 202648
rect 323032 202700 323084 202706
rect 323032 202642 323084 202648
rect 333900 202638 333928 205006
rect 344296 202638 344324 226306
rect 345018 214568 345074 214577
rect 345018 214503 345074 214512
rect 345032 205562 345060 214503
rect 345020 205556 345072 205562
rect 345020 205498 345072 205504
rect 345676 205494 345704 226442
rect 352012 226432 352064 226438
rect 352012 226374 352064 226380
rect 352024 224876 352052 226374
rect 361684 224876 361712 226442
rect 371332 226364 371384 226370
rect 371332 226306 371384 226312
rect 371344 224876 371372 226306
rect 350446 215248 350502 215257
rect 350446 215183 350502 215192
rect 350460 205562 350488 215183
rect 371528 205714 371556 226442
rect 374644 226432 374696 226438
rect 374644 226374 374696 226380
rect 373264 226364 373316 226370
rect 373264 226306 373316 226312
rect 371358 205686 371556 205714
rect 350448 205556 350500 205562
rect 350448 205498 350500 205504
rect 345664 205488 345716 205494
rect 345664 205430 345716 205436
rect 352024 202706 352052 205020
rect 361684 202706 361712 205020
rect 373276 202706 373304 226306
rect 373998 214568 374054 214577
rect 373998 214503 374054 214512
rect 374012 205630 374040 214503
rect 374000 205624 374052 205630
rect 374000 205566 374052 205572
rect 374656 202842 374684 226374
rect 389376 224890 389404 226442
rect 399024 226364 399076 226370
rect 399024 226306 399076 226312
rect 399036 224890 399064 226306
rect 389376 224862 389712 224890
rect 399036 224862 399372 224890
rect 379624 224318 380052 224346
rect 378046 215248 378102 215257
rect 378046 215183 378102 215192
rect 378060 205494 378088 215183
rect 378048 205488 378100 205494
rect 378048 205430 378100 205436
rect 374644 202836 374696 202842
rect 374644 202778 374696 202784
rect 379624 202706 379652 224318
rect 399496 205714 399524 226442
rect 400864 226364 400916 226370
rect 400864 226306 400916 226312
rect 399372 205686 399524 205714
rect 379716 205006 380052 205034
rect 389712 205006 390048 205034
rect 379716 202842 379744 205006
rect 379704 202836 379756 202842
rect 379704 202778 379756 202784
rect 352012 202700 352064 202706
rect 352012 202642 352064 202648
rect 361672 202700 361724 202706
rect 361672 202642 361724 202648
rect 373264 202700 373316 202706
rect 373264 202642 373316 202648
rect 379612 202700 379664 202706
rect 379612 202642 379664 202648
rect 390020 202638 390048 205006
rect 400876 202638 400904 226306
rect 408052 224876 408080 226510
rect 417700 226500 417752 226506
rect 417700 226442 417752 226448
rect 417712 224876 417740 226442
rect 428556 226432 428608 226438
rect 428556 226374 428608 226380
rect 427360 226364 427412 226370
rect 427360 226306 427412 226312
rect 428464 226364 428516 226370
rect 428464 226306 428516 226312
rect 427372 224876 427400 226306
rect 405646 215248 405702 215257
rect 405646 215183 405702 215192
rect 401598 214568 401654 214577
rect 401598 214503 401654 214512
rect 401612 205562 401640 214503
rect 405660 205630 405688 215183
rect 405648 205624 405700 205630
rect 405648 205566 405700 205572
rect 427386 205562 427768 205578
rect 401600 205556 401652 205562
rect 427386 205556 427780 205562
rect 427386 205550 427728 205556
rect 401600 205498 401652 205504
rect 427728 205498 427780 205504
rect 408052 202706 408080 205020
rect 417712 202706 417740 205020
rect 428476 202706 428504 226306
rect 428568 205562 428596 226374
rect 428660 207670 428688 226510
rect 456156 226500 456208 226506
rect 456156 226442 456208 226448
rect 473360 226500 473412 226506
rect 473360 226442 473412 226448
rect 483480 226500 483532 226506
rect 483480 226442 483532 226448
rect 445668 226432 445720 226438
rect 445668 226374 445720 226380
rect 445680 224876 445708 226374
rect 455328 226364 455380 226370
rect 455328 226306 455380 226312
rect 456064 226364 456116 226370
rect 456064 226306 456116 226312
rect 455340 224876 455368 226306
rect 434824 224318 436034 224346
rect 434626 215248 434682 215257
rect 434626 215183 434682 215192
rect 429198 214568 429254 214577
rect 429198 214503 429254 214512
rect 428648 207664 428700 207670
rect 428648 207606 428700 207612
rect 428556 205556 428608 205562
rect 428556 205498 428608 205504
rect 429212 205494 429240 214503
rect 434640 205562 434668 215183
rect 434628 205556 434680 205562
rect 434628 205498 434680 205504
rect 429200 205488 429252 205494
rect 429200 205430 429252 205436
rect 434824 202706 434852 224318
rect 435732 207664 435784 207670
rect 435732 207606 435784 207612
rect 435744 205714 435772 207606
rect 455696 207392 455748 207398
rect 455696 207334 455748 207340
rect 455708 205714 455736 207334
rect 435744 205686 436034 205714
rect 455354 205686 455736 205714
rect 408040 202700 408092 202706
rect 408040 202642 408092 202648
rect 417700 202700 417752 202706
rect 417700 202642 417752 202648
rect 428464 202700 428516 202706
rect 428464 202642 428516 202648
rect 434812 202700 434864 202706
rect 434812 202642 434864 202648
rect 445680 202638 445708 205020
rect 456076 202638 456104 226306
rect 456168 207398 456196 226442
rect 464344 226432 464396 226438
rect 464344 226374 464396 226380
rect 464356 224890 464384 226374
rect 464048 224862 464384 224890
rect 473372 224890 473400 226442
rect 483020 226364 483072 226370
rect 483020 226306 483072 226312
rect 483032 224890 483060 226306
rect 473372 224862 473708 224890
rect 483032 224862 483368 224890
rect 462226 215248 462282 215257
rect 462226 215183 462282 215192
rect 458178 214568 458234 214577
rect 458178 214503 458234 214512
rect 456156 207392 456208 207398
rect 456156 207334 456208 207340
rect 458192 205630 458220 214503
rect 458180 205624 458232 205630
rect 458180 205566 458232 205572
rect 462240 205494 462268 215183
rect 483492 205714 483520 226442
rect 483664 226432 483716 226438
rect 483664 226374 483716 226380
rect 483676 207466 483704 226374
rect 485044 226364 485096 226370
rect 485044 226306 485096 226312
rect 483664 207460 483716 207466
rect 483664 207402 483716 207408
rect 483368 205686 483520 205714
rect 462228 205488 462280 205494
rect 462228 205430 462280 205436
rect 463712 205006 464048 205034
rect 473708 205006 474044 205034
rect 463712 202706 463740 205006
rect 474016 202706 474044 205006
rect 485056 202706 485084 226306
rect 489826 215248 489882 215257
rect 489826 215183 489882 215192
rect 485778 214568 485834 214577
rect 485778 214503 485834 214512
rect 485792 205562 485820 214503
rect 489840 205630 489868 215183
rect 489828 205624 489880 205630
rect 489828 205566 489880 205572
rect 485780 205556 485832 205562
rect 485780 205498 485832 205504
rect 463700 202700 463752 202706
rect 463700 202642 463752 202648
rect 474004 202700 474056 202706
rect 474004 202642 474056 202648
rect 485044 202700 485096 202706
rect 485044 202642 485096 202648
rect 333888 202632 333940 202638
rect 333888 202574 333940 202580
rect 344284 202632 344336 202638
rect 344284 202574 344336 202580
rect 390008 202632 390060 202638
rect 390008 202574 390060 202580
rect 400864 202632 400916 202638
rect 400864 202574 400916 202580
rect 445668 202632 445720 202638
rect 445668 202574 445720 202580
rect 456064 202632 456116 202638
rect 456064 202574 456116 202580
rect 296352 200388 296404 200394
rect 296352 200330 296404 200336
rect 316776 200388 316828 200394
rect 316776 200330 316828 200336
rect 408040 200388 408092 200394
rect 408040 200330 408092 200336
rect 428648 200388 428700 200394
rect 428648 200330 428700 200336
rect 277676 200320 277728 200326
rect 277676 200262 277728 200268
rect 287520 200320 287572 200326
rect 287520 200262 287572 200268
rect 268016 200252 268068 200258
rect 268016 200194 268068 200200
rect 268028 197948 268056 200194
rect 277688 197948 277716 200262
rect 287336 200184 287388 200190
rect 287336 200126 287388 200132
rect 287348 197948 287376 200126
rect 266266 188320 266322 188329
rect 266266 188255 266322 188264
rect 262218 187640 262274 187649
rect 262218 187575 262274 187584
rect 262232 179382 262260 187575
rect 266280 179382 266308 188255
rect 262220 179376 262272 179382
rect 262220 179318 262272 179324
rect 266268 179376 266320 179382
rect 266268 179318 266320 179324
rect 287532 178786 287560 200262
rect 287704 200252 287756 200258
rect 287704 200194 287756 200200
rect 287716 179450 287744 200194
rect 289084 200184 289136 200190
rect 289084 200126 289136 200132
rect 287704 179444 287756 179450
rect 287704 179386 287756 179392
rect 287362 178758 287560 178786
rect 249708 176588 249760 176594
rect 249708 176530 249760 176536
rect 260104 176588 260156 176594
rect 260104 176530 260156 176536
rect 261484 176588 261536 176594
rect 261484 176530 261536 176536
rect 268028 176526 268056 178092
rect 277688 176526 277716 178092
rect 289096 176526 289124 200126
rect 296364 197962 296392 200330
rect 305368 200320 305420 200326
rect 305368 200262 305420 200268
rect 296056 197934 296392 197962
rect 305380 197962 305408 200262
rect 315488 200252 315540 200258
rect 315488 200194 315540 200200
rect 315028 200184 315080 200190
rect 315028 200126 315080 200132
rect 315040 197962 315068 200126
rect 305380 197934 305716 197962
rect 315040 197934 315376 197962
rect 293866 188320 293922 188329
rect 293866 188255 293922 188264
rect 289818 187640 289874 187649
rect 289818 187575 289874 187584
rect 289832 179314 289860 187575
rect 293880 179314 293908 188255
rect 295708 179444 295760 179450
rect 295708 179386 295760 179392
rect 289820 179308 289872 179314
rect 289820 179250 289872 179256
rect 293868 179308 293920 179314
rect 293868 179250 293920 179256
rect 295720 178786 295748 179386
rect 315500 178786 315528 200194
rect 316684 200184 316736 200190
rect 316684 200126 316736 200132
rect 295720 178758 296056 178786
rect 315376 178758 315528 178786
rect 305716 178078 306052 178106
rect 306024 176526 306052 178078
rect 316696 176526 316724 200126
rect 316788 179450 316816 200330
rect 345664 200320 345716 200326
rect 345664 200262 345716 200268
rect 361672 200320 361724 200326
rect 361672 200262 361724 200268
rect 371516 200320 371568 200326
rect 371516 200262 371568 200268
rect 389364 200320 389416 200326
rect 389364 200262 389416 200268
rect 399484 200320 399536 200326
rect 399484 200262 399536 200268
rect 333704 200252 333756 200258
rect 333704 200194 333756 200200
rect 333716 197948 333744 200194
rect 343364 200184 343416 200190
rect 343364 200126 343416 200132
rect 344284 200184 344336 200190
rect 344284 200126 344336 200132
rect 343376 197948 343404 200126
rect 323044 197254 324070 197282
rect 322846 188320 322902 188329
rect 322846 188255 322902 188264
rect 317418 187640 317474 187649
rect 317418 187575 317474 187584
rect 316776 179444 316828 179450
rect 316776 179386 316828 179392
rect 317432 179382 317460 187575
rect 322860 179382 322888 188255
rect 317420 179376 317472 179382
rect 317420 179318 317472 179324
rect 322848 179376 322900 179382
rect 322848 179318 322900 179324
rect 323044 176526 323072 197254
rect 323676 179444 323728 179450
rect 323676 179386 323728 179392
rect 323688 178786 323716 179386
rect 343548 179308 343600 179314
rect 343548 179250 343600 179256
rect 343560 178786 343588 179250
rect 323688 178758 324070 178786
rect 343390 178758 343588 178786
rect 238852 176520 238904 176526
rect 238852 176462 238904 176468
rect 268016 176520 268068 176526
rect 268016 176462 268068 176468
rect 277676 176520 277728 176526
rect 277676 176462 277728 176468
rect 289084 176520 289136 176526
rect 289084 176462 289136 176468
rect 306012 176520 306064 176526
rect 306012 176462 306064 176468
rect 316684 176520 316736 176526
rect 316684 176462 316736 176468
rect 323032 176520 323084 176526
rect 323032 176462 323084 176468
rect 333716 176458 333744 178092
rect 344296 176458 344324 200126
rect 345018 187640 345074 187649
rect 345018 187575 345074 187584
rect 345032 179246 345060 187575
rect 345676 179314 345704 200262
rect 352012 200252 352064 200258
rect 352012 200194 352064 200200
rect 352024 197948 352052 200194
rect 361684 197948 361712 200262
rect 371332 200184 371384 200190
rect 371332 200126 371384 200132
rect 371344 197948 371372 200126
rect 350446 188320 350502 188329
rect 350446 188255 350502 188264
rect 350460 179314 350488 188255
rect 345664 179308 345716 179314
rect 345664 179250 345716 179256
rect 350448 179308 350500 179314
rect 350448 179250 350500 179256
rect 345020 179240 345072 179246
rect 345020 179182 345072 179188
rect 371528 178786 371556 200262
rect 374644 200252 374696 200258
rect 374644 200194 374696 200200
rect 373264 200184 373316 200190
rect 373264 200126 373316 200132
rect 371358 178758 371556 178786
rect 352024 176526 352052 178092
rect 361684 176526 361712 178092
rect 373276 176526 373304 200126
rect 373998 187640 374054 187649
rect 373998 187575 374054 187584
rect 374012 179382 374040 187575
rect 374000 179376 374052 179382
rect 374000 179318 374052 179324
rect 374656 176662 374684 200194
rect 389376 197962 389404 200262
rect 399024 200184 399076 200190
rect 399024 200126 399076 200132
rect 399036 197962 399064 200126
rect 389376 197934 389712 197962
rect 399036 197934 399372 197962
rect 379624 197254 380052 197282
rect 378046 188320 378102 188329
rect 378046 188255 378102 188264
rect 378060 179246 378088 188255
rect 378048 179240 378100 179246
rect 378048 179182 378100 179188
rect 374644 176656 374696 176662
rect 374644 176598 374696 176604
rect 379624 176526 379652 197254
rect 399496 178786 399524 200262
rect 400864 200184 400916 200190
rect 400864 200126 400916 200132
rect 399372 178758 399524 178786
rect 379716 178078 380052 178106
rect 389712 178078 390048 178106
rect 379716 176662 379744 178078
rect 379704 176656 379756 176662
rect 379704 176598 379756 176604
rect 352012 176520 352064 176526
rect 352012 176462 352064 176468
rect 361672 176520 361724 176526
rect 361672 176462 361724 176468
rect 373264 176520 373316 176526
rect 373264 176462 373316 176468
rect 379612 176520 379664 176526
rect 379612 176462 379664 176468
rect 390020 176458 390048 178078
rect 400876 176458 400904 200126
rect 408052 197948 408080 200330
rect 417700 200320 417752 200326
rect 417700 200262 417752 200268
rect 417712 197948 417740 200262
rect 428464 200252 428516 200258
rect 428464 200194 428516 200200
rect 427360 200184 427412 200190
rect 427360 200126 427412 200132
rect 427372 197948 427400 200126
rect 405646 188320 405702 188329
rect 405646 188255 405702 188264
rect 401598 187640 401654 187649
rect 401598 187575 401654 187584
rect 401612 179314 401640 187575
rect 405660 179382 405688 188255
rect 428476 180794 428504 200194
rect 428556 200184 428608 200190
rect 428556 200126 428608 200132
rect 427832 180766 428504 180794
rect 405648 179376 405700 179382
rect 405648 179318 405700 179324
rect 401600 179308 401652 179314
rect 401600 179250 401652 179256
rect 427832 178786 427860 180766
rect 427386 178758 427860 178786
rect 408052 176526 408080 178092
rect 417712 176526 417740 178092
rect 428568 176526 428596 200126
rect 428660 180130 428688 200330
rect 456156 200320 456208 200326
rect 456156 200262 456208 200268
rect 473544 200320 473596 200326
rect 473544 200262 473596 200268
rect 483480 200320 483532 200326
rect 483480 200262 483532 200268
rect 445668 200252 445720 200258
rect 445668 200194 445720 200200
rect 445680 197948 445708 200194
rect 455328 200184 455380 200190
rect 455328 200126 455380 200132
rect 456064 200184 456116 200190
rect 456064 200126 456116 200132
rect 455340 197948 455368 200126
rect 434824 197254 436034 197282
rect 434626 188320 434682 188329
rect 434626 188255 434682 188264
rect 429198 187640 429254 187649
rect 429198 187575 429254 187584
rect 428648 180124 428700 180130
rect 428648 180066 428700 180072
rect 429212 179246 429240 187575
rect 434640 179314 434668 188255
rect 434628 179308 434680 179314
rect 434628 179250 434680 179256
rect 429200 179240 429252 179246
rect 429200 179182 429252 179188
rect 434824 176526 434852 197254
rect 455696 185632 455748 185638
rect 455696 185574 455748 185580
rect 435732 180124 435784 180130
rect 435732 180066 435784 180072
rect 435744 178786 435772 180066
rect 455708 178786 455736 185574
rect 435744 178758 436034 178786
rect 455354 178758 455736 178786
rect 408040 176520 408092 176526
rect 408040 176462 408092 176468
rect 417700 176520 417752 176526
rect 417700 176462 417752 176468
rect 428556 176520 428608 176526
rect 428556 176462 428608 176468
rect 434812 176520 434864 176526
rect 434812 176462 434864 176468
rect 445680 176458 445708 178092
rect 456076 176458 456104 200126
rect 456168 185638 456196 200262
rect 464344 200252 464396 200258
rect 464344 200194 464396 200200
rect 464356 197962 464384 200194
rect 464048 197934 464384 197962
rect 473556 197962 473584 200262
rect 483204 200184 483256 200190
rect 483204 200126 483256 200132
rect 483216 197962 483244 200126
rect 473556 197934 473708 197962
rect 483216 197934 483368 197962
rect 462226 188320 462282 188329
rect 462226 188255 462282 188264
rect 458178 187640 458234 187649
rect 458178 187575 458234 187584
rect 456156 185632 456208 185638
rect 456156 185574 456208 185580
rect 458192 179382 458220 187575
rect 458180 179376 458232 179382
rect 458180 179318 458232 179324
rect 462240 179246 462268 188255
rect 462228 179240 462280 179246
rect 462228 179182 462280 179188
rect 483492 178786 483520 200262
rect 483664 200252 483716 200258
rect 483664 200194 483716 200200
rect 483676 179722 483704 200194
rect 485044 200184 485096 200190
rect 485044 200126 485096 200132
rect 483664 179716 483716 179722
rect 483664 179658 483716 179664
rect 483368 178758 483520 178786
rect 463712 178078 464048 178106
rect 473708 178078 474044 178106
rect 463712 176526 463740 178078
rect 474016 176526 474044 178078
rect 485056 176526 485084 200126
rect 489826 188320 489882 188329
rect 489826 188255 489882 188264
rect 485778 187640 485834 187649
rect 485778 187575 485834 187584
rect 485792 179314 485820 187575
rect 489840 179382 489868 188255
rect 489828 179376 489880 179382
rect 489828 179318 489880 179324
rect 485780 179308 485832 179314
rect 485780 179250 485832 179256
rect 463700 176520 463752 176526
rect 463700 176462 463752 176468
rect 474004 176520 474056 176526
rect 474004 176462 474056 176468
rect 485044 176520 485096 176526
rect 485044 176462 485096 176468
rect 333704 176452 333756 176458
rect 333704 176394 333756 176400
rect 344284 176452 344336 176458
rect 344284 176394 344336 176400
rect 390008 176452 390060 176458
rect 390008 176394 390060 176400
rect 400864 176452 400916 176458
rect 400864 176394 400916 176400
rect 445668 176452 445720 176458
rect 445668 176394 445720 176400
rect 456064 176452 456116 176458
rect 456064 176394 456116 176400
rect 296352 172780 296404 172786
rect 296352 172722 296404 172728
rect 316776 172780 316828 172786
rect 316776 172722 316828 172728
rect 408040 172780 408092 172786
rect 408040 172722 408092 172728
rect 428648 172780 428700 172786
rect 428648 172722 428700 172728
rect 260196 172712 260248 172718
rect 260196 172654 260248 172660
rect 277676 172712 277728 172718
rect 277676 172654 277728 172660
rect 287520 172712 287572 172718
rect 287520 172654 287572 172660
rect 249708 172644 249760 172650
rect 249708 172586 249760 172592
rect 249720 170884 249748 172586
rect 259368 172576 259420 172582
rect 259368 172518 259420 172524
rect 260104 172576 260156 172582
rect 260104 172518 260156 172524
rect 259380 170884 259408 172518
rect 238864 170326 240074 170354
rect 238666 161256 238722 161265
rect 238666 161191 238722 161200
rect 238680 151706 238708 161191
rect 238668 151700 238720 151706
rect 238668 151642 238720 151648
rect 238864 148918 238892 170326
rect 259736 156664 259788 156670
rect 259736 156606 259788 156612
rect 239772 152584 239824 152590
rect 239772 152526 239824 152532
rect 239784 151722 239812 152526
rect 259748 151722 259776 156606
rect 239784 151694 240074 151722
rect 259394 151694 259776 151722
rect 238852 148912 238904 148918
rect 238852 148854 238904 148860
rect 249720 148850 249748 151028
rect 260116 148850 260144 172518
rect 260208 156670 260236 172654
rect 268016 172644 268068 172650
rect 268016 172586 268068 172592
rect 268028 170884 268056 172586
rect 277688 170884 277716 172654
rect 287336 172576 287388 172582
rect 287336 172518 287388 172524
rect 287348 170884 287376 172518
rect 266266 161256 266322 161265
rect 266266 161191 266322 161200
rect 262218 160576 262274 160585
rect 262218 160511 262274 160520
rect 260196 156664 260248 156670
rect 260196 156606 260248 156612
rect 262232 151774 262260 160511
rect 266280 151774 266308 161191
rect 262220 151768 262272 151774
rect 262220 151710 262272 151716
rect 266268 151768 266320 151774
rect 287532 151722 287560 172654
rect 287704 172644 287756 172650
rect 287704 172586 287756 172592
rect 287716 153202 287744 172586
rect 289084 172576 289136 172582
rect 289084 172518 289136 172524
rect 287704 153196 287756 153202
rect 287704 153138 287756 153144
rect 266268 151710 266320 151716
rect 287362 151694 287560 151722
rect 268028 148918 268056 151028
rect 277688 148918 277716 151028
rect 289096 148918 289124 172518
rect 296364 170898 296392 172722
rect 305368 172712 305420 172718
rect 305368 172654 305420 172660
rect 296056 170870 296392 170898
rect 305380 170898 305408 172654
rect 315488 172644 315540 172650
rect 315488 172586 315540 172592
rect 315028 172576 315080 172582
rect 315028 172518 315080 172524
rect 315040 170898 315068 172518
rect 305380 170870 305716 170898
rect 315040 170870 315376 170898
rect 293866 161256 293922 161265
rect 293866 161191 293922 161200
rect 289818 160576 289874 160585
rect 289818 160511 289874 160520
rect 289832 151706 289860 160511
rect 293880 151706 293908 161191
rect 295708 153196 295760 153202
rect 295708 153138 295760 153144
rect 295720 151722 295748 153138
rect 315500 151722 315528 172586
rect 316684 172576 316736 172582
rect 316684 172518 316736 172524
rect 289820 151700 289872 151706
rect 289820 151642 289872 151648
rect 293868 151700 293920 151706
rect 295720 151694 296056 151722
rect 315376 151694 315528 151722
rect 293868 151642 293920 151648
rect 305716 151014 306052 151042
rect 306024 148918 306052 151014
rect 316696 148918 316724 172518
rect 316788 153202 316816 172722
rect 345664 172712 345716 172718
rect 345664 172654 345716 172660
rect 361672 172712 361724 172718
rect 361672 172654 361724 172660
rect 371516 172712 371568 172718
rect 371516 172654 371568 172660
rect 389364 172712 389416 172718
rect 389364 172654 389416 172660
rect 399484 172712 399536 172718
rect 399484 172654 399536 172660
rect 333704 172644 333756 172650
rect 333704 172586 333756 172592
rect 333716 170884 333744 172586
rect 343364 172576 343416 172582
rect 343364 172518 343416 172524
rect 344284 172576 344336 172582
rect 344284 172518 344336 172524
rect 343376 170884 343404 172518
rect 323044 170326 324070 170354
rect 322846 161256 322902 161265
rect 322846 161191 322902 161200
rect 317418 160576 317474 160585
rect 317418 160511 317474 160520
rect 316776 153196 316828 153202
rect 316776 153138 316828 153144
rect 317432 151774 317460 160511
rect 322860 151774 322888 161191
rect 317420 151768 317472 151774
rect 317420 151710 317472 151716
rect 322848 151768 322900 151774
rect 322848 151710 322900 151716
rect 323044 148918 323072 170326
rect 323676 153196 323728 153202
rect 323676 153138 323728 153144
rect 323688 151722 323716 153138
rect 323688 151694 324070 151722
rect 343390 151706 343680 151722
rect 343390 151700 343692 151706
rect 343390 151694 343640 151700
rect 343640 151642 343692 151648
rect 268016 148912 268068 148918
rect 268016 148854 268068 148860
rect 277676 148912 277728 148918
rect 277676 148854 277728 148860
rect 289084 148912 289136 148918
rect 289084 148854 289136 148860
rect 306012 148912 306064 148918
rect 306012 148854 306064 148860
rect 316684 148912 316736 148918
rect 316684 148854 316736 148860
rect 323032 148912 323084 148918
rect 323032 148854 323084 148860
rect 333716 148850 333744 151028
rect 344296 148850 344324 172518
rect 345018 160576 345074 160585
rect 345018 160511 345074 160520
rect 345032 151638 345060 160511
rect 345676 151706 345704 172654
rect 352012 172644 352064 172650
rect 352012 172586 352064 172592
rect 352024 170884 352052 172586
rect 361684 170884 361712 172654
rect 371332 172576 371384 172582
rect 371332 172518 371384 172524
rect 371344 170884 371372 172518
rect 350446 161256 350502 161265
rect 350446 161191 350502 161200
rect 350460 151706 350488 161191
rect 371528 151722 371556 172654
rect 374644 172644 374696 172650
rect 374644 172586 374696 172592
rect 373264 172576 373316 172582
rect 373264 172518 373316 172524
rect 345664 151700 345716 151706
rect 345664 151642 345716 151648
rect 350448 151700 350500 151706
rect 371358 151694 371556 151722
rect 350448 151642 350500 151648
rect 345020 151632 345072 151638
rect 345020 151574 345072 151580
rect 352024 148918 352052 151028
rect 361684 148918 361712 151028
rect 373276 148918 373304 172518
rect 373998 160576 374054 160585
rect 373998 160511 374054 160520
rect 374012 151774 374040 160511
rect 374000 151768 374052 151774
rect 374000 151710 374052 151716
rect 374656 149054 374684 172586
rect 389376 170898 389404 172654
rect 399024 172576 399076 172582
rect 399024 172518 399076 172524
rect 399036 170898 399064 172518
rect 389376 170870 389712 170898
rect 399036 170870 399372 170898
rect 379624 170326 380052 170354
rect 378046 161256 378102 161265
rect 378046 161191 378102 161200
rect 378060 151638 378088 161191
rect 378048 151632 378100 151638
rect 378048 151574 378100 151580
rect 374644 149048 374696 149054
rect 374644 148990 374696 148996
rect 379624 148918 379652 170326
rect 399496 151722 399524 172654
rect 400864 172576 400916 172582
rect 400864 172518 400916 172524
rect 399372 151694 399524 151722
rect 379716 151014 380052 151042
rect 389712 151014 390048 151042
rect 379716 149054 379744 151014
rect 379704 149048 379756 149054
rect 379704 148990 379756 148996
rect 352012 148912 352064 148918
rect 352012 148854 352064 148860
rect 361672 148912 361724 148918
rect 361672 148854 361724 148860
rect 373264 148912 373316 148918
rect 373264 148854 373316 148860
rect 379612 148912 379664 148918
rect 379612 148854 379664 148860
rect 390020 148850 390048 151014
rect 400876 148850 400904 172518
rect 408052 170884 408080 172722
rect 417700 172712 417752 172718
rect 417700 172654 417752 172660
rect 417712 170884 417740 172654
rect 428464 172644 428516 172650
rect 428464 172586 428516 172592
rect 427360 172576 427412 172582
rect 427360 172518 427412 172524
rect 427372 170884 427400 172518
rect 405646 161256 405702 161265
rect 405646 161191 405702 161200
rect 401598 160576 401654 160585
rect 401598 160511 401654 160520
rect 401612 151706 401640 160511
rect 405660 151774 405688 161191
rect 428476 151814 428504 172586
rect 428556 172576 428608 172582
rect 428556 172518 428608 172524
rect 427832 151786 428504 151814
rect 405648 151768 405700 151774
rect 427832 151722 427860 151786
rect 405648 151710 405700 151716
rect 401600 151700 401652 151706
rect 427386 151694 427860 151722
rect 401600 151642 401652 151648
rect 408052 148918 408080 151028
rect 417712 148918 417740 151028
rect 428568 148918 428596 172518
rect 428660 152522 428688 172722
rect 456156 172712 456208 172718
rect 456156 172654 456208 172660
rect 473544 172712 473596 172718
rect 473544 172654 473596 172660
rect 483480 172712 483532 172718
rect 483480 172654 483532 172660
rect 445668 172644 445720 172650
rect 445668 172586 445720 172592
rect 445680 170884 445708 172586
rect 455328 172576 455380 172582
rect 455328 172518 455380 172524
rect 456064 172576 456116 172582
rect 456064 172518 456116 172524
rect 455340 170884 455368 172518
rect 434824 170326 436034 170354
rect 434626 161256 434682 161265
rect 434626 161191 434682 161200
rect 429198 160576 429254 160585
rect 429198 160511 429254 160520
rect 428648 152516 428700 152522
rect 428648 152458 428700 152464
rect 429212 151638 429240 160511
rect 434640 151706 434668 161191
rect 434628 151700 434680 151706
rect 434628 151642 434680 151648
rect 429200 151632 429252 151638
rect 429200 151574 429252 151580
rect 434824 148918 434852 170326
rect 455696 156664 455748 156670
rect 455696 156606 455748 156612
rect 435732 152516 435784 152522
rect 435732 152458 435784 152464
rect 435744 151722 435772 152458
rect 455708 151722 455736 156606
rect 435744 151694 436034 151722
rect 455354 151694 455736 151722
rect 408040 148912 408092 148918
rect 408040 148854 408092 148860
rect 417700 148912 417752 148918
rect 417700 148854 417752 148860
rect 428556 148912 428608 148918
rect 428556 148854 428608 148860
rect 434812 148912 434864 148918
rect 434812 148854 434864 148860
rect 445680 148850 445708 151028
rect 456076 148850 456104 172518
rect 456168 156670 456196 172654
rect 464344 172644 464396 172650
rect 464344 172586 464396 172592
rect 464356 170898 464384 172586
rect 464048 170870 464384 170898
rect 473556 170898 473584 172654
rect 483204 172576 483256 172582
rect 483204 172518 483256 172524
rect 483216 170898 483244 172518
rect 473556 170870 473708 170898
rect 483216 170870 483368 170898
rect 462226 161256 462282 161265
rect 462226 161191 462282 161200
rect 458178 160576 458234 160585
rect 458178 160511 458234 160520
rect 456156 156664 456208 156670
rect 456156 156606 456208 156612
rect 458192 151774 458220 160511
rect 458180 151768 458232 151774
rect 458180 151710 458232 151716
rect 462240 151638 462268 161191
rect 483492 151722 483520 172654
rect 483664 172644 483716 172650
rect 483664 172586 483716 172592
rect 483676 152522 483704 172586
rect 485044 172576 485096 172582
rect 485044 172518 485096 172524
rect 483664 152516 483716 152522
rect 483664 152458 483716 152464
rect 483368 151694 483520 151722
rect 462228 151632 462280 151638
rect 462228 151574 462280 151580
rect 463712 151014 464048 151042
rect 473708 151014 474044 151042
rect 463712 148918 463740 151014
rect 474016 148918 474044 151014
rect 485056 148918 485084 172518
rect 489826 161256 489882 161265
rect 489826 161191 489882 161200
rect 485778 160576 485834 160585
rect 485778 160511 485834 160520
rect 485792 151706 485820 160511
rect 489840 151774 489868 161191
rect 489828 151768 489880 151774
rect 489828 151710 489880 151716
rect 485780 151700 485832 151706
rect 485780 151642 485832 151648
rect 463700 148912 463752 148918
rect 463700 148854 463752 148860
rect 474004 148912 474056 148918
rect 474004 148854 474056 148860
rect 485044 148912 485096 148918
rect 485044 148854 485096 148860
rect 249708 148844 249760 148850
rect 249708 148786 249760 148792
rect 260104 148844 260156 148850
rect 260104 148786 260156 148792
rect 333704 148844 333756 148850
rect 333704 148786 333756 148792
rect 344284 148844 344336 148850
rect 344284 148786 344336 148792
rect 390008 148844 390060 148850
rect 390008 148786 390060 148792
rect 400864 148844 400916 148850
rect 400864 148786 400916 148792
rect 445668 148844 445720 148850
rect 445668 148786 445720 148792
rect 456064 148844 456116 148850
rect 456064 148786 456116 148792
rect 296352 146532 296404 146538
rect 296352 146474 296404 146480
rect 316776 146532 316828 146538
rect 316776 146474 316828 146480
rect 408040 146532 408092 146538
rect 408040 146474 408092 146480
rect 428648 146532 428700 146538
rect 428648 146474 428700 146480
rect 260104 146464 260156 146470
rect 260104 146406 260156 146412
rect 277676 146464 277728 146470
rect 277676 146406 277728 146412
rect 287520 146464 287572 146470
rect 287520 146406 287572 146412
rect 249708 146396 249760 146402
rect 249708 146338 249760 146344
rect 249720 143956 249748 146338
rect 259368 146328 259420 146334
rect 259368 146270 259420 146276
rect 259380 143956 259408 146270
rect 238864 143262 240074 143290
rect 238666 134328 238722 134337
rect 238666 134263 238722 134272
rect 238680 125526 238708 134263
rect 238668 125520 238720 125526
rect 238668 125462 238720 125468
rect 238864 122670 238892 143262
rect 260116 132494 260144 146406
rect 268016 146396 268068 146402
rect 268016 146338 268068 146344
rect 260196 146328 260248 146334
rect 260196 146270 260248 146276
rect 259840 132466 260144 132494
rect 239772 126948 239824 126954
rect 239772 126890 239824 126896
rect 239784 124794 239812 126890
rect 259840 124794 259868 132466
rect 239784 124766 240074 124794
rect 259394 124766 259868 124794
rect 238852 122664 238904 122670
rect 238852 122606 238904 122612
rect 249720 122602 249748 124100
rect 260208 122602 260236 146270
rect 268028 143956 268056 146338
rect 277688 143956 277716 146406
rect 287336 146328 287388 146334
rect 287336 146270 287388 146276
rect 287348 143956 287376 146270
rect 266266 134328 266322 134337
rect 266266 134263 266322 134272
rect 262218 133648 262274 133657
rect 262218 133583 262274 133592
rect 262232 125594 262260 133583
rect 266280 125594 266308 134263
rect 262220 125588 262272 125594
rect 262220 125530 262272 125536
rect 266268 125588 266320 125594
rect 266268 125530 266320 125536
rect 287532 124794 287560 146406
rect 287704 146396 287756 146402
rect 287704 146338 287756 146344
rect 287716 126138 287744 146338
rect 289084 146328 289136 146334
rect 289084 146270 289136 146276
rect 287704 126132 287756 126138
rect 287704 126074 287756 126080
rect 287362 124766 287560 124794
rect 268028 122670 268056 124100
rect 277688 122670 277716 124100
rect 289096 122670 289124 146270
rect 296364 143970 296392 146474
rect 305368 146464 305420 146470
rect 305368 146406 305420 146412
rect 296056 143942 296392 143970
rect 305380 143970 305408 146406
rect 315488 146396 315540 146402
rect 315488 146338 315540 146344
rect 315028 146328 315080 146334
rect 315028 146270 315080 146276
rect 315040 143970 315068 146270
rect 305380 143942 305716 143970
rect 315040 143942 315376 143970
rect 293866 134328 293922 134337
rect 293866 134263 293922 134272
rect 289818 133648 289874 133657
rect 289818 133583 289874 133592
rect 289832 125526 289860 133583
rect 293880 125526 293908 134263
rect 295708 126132 295760 126138
rect 295708 126074 295760 126080
rect 289820 125520 289872 125526
rect 289820 125462 289872 125468
rect 293868 125520 293920 125526
rect 293868 125462 293920 125468
rect 295720 124794 295748 126074
rect 315500 124794 315528 146338
rect 316684 146328 316736 146334
rect 316684 146270 316736 146276
rect 295720 124766 296056 124794
rect 315376 124766 315528 124794
rect 305716 124086 306052 124114
rect 306024 122670 306052 124086
rect 316696 122670 316724 146270
rect 316788 126138 316816 146474
rect 345664 146464 345716 146470
rect 345664 146406 345716 146412
rect 361672 146464 361724 146470
rect 361672 146406 361724 146412
rect 371516 146464 371568 146470
rect 371516 146406 371568 146412
rect 389364 146464 389416 146470
rect 389364 146406 389416 146412
rect 399484 146464 399536 146470
rect 399484 146406 399536 146412
rect 333704 146396 333756 146402
rect 333704 146338 333756 146344
rect 333716 143956 333744 146338
rect 343364 146328 343416 146334
rect 343364 146270 343416 146276
rect 344284 146328 344336 146334
rect 344284 146270 344336 146276
rect 343376 143956 343404 146270
rect 323044 143262 324070 143290
rect 322846 134328 322902 134337
rect 322846 134263 322902 134272
rect 317418 133648 317474 133657
rect 317418 133583 317474 133592
rect 316776 126132 316828 126138
rect 316776 126074 316828 126080
rect 317432 125594 317460 133583
rect 322860 125594 322888 134263
rect 317420 125588 317472 125594
rect 317420 125530 317472 125536
rect 322848 125588 322900 125594
rect 322848 125530 322900 125536
rect 323044 122670 323072 143262
rect 323676 126132 323728 126138
rect 323676 126074 323728 126080
rect 323688 124794 323716 126074
rect 343548 124840 343600 124846
rect 323688 124766 324070 124794
rect 343390 124788 343548 124794
rect 343390 124782 343600 124788
rect 343390 124766 343588 124782
rect 268016 122664 268068 122670
rect 268016 122606 268068 122612
rect 277676 122664 277728 122670
rect 277676 122606 277728 122612
rect 289084 122664 289136 122670
rect 289084 122606 289136 122612
rect 306012 122664 306064 122670
rect 306012 122606 306064 122612
rect 316684 122664 316736 122670
rect 316684 122606 316736 122612
rect 323032 122664 323084 122670
rect 323032 122606 323084 122612
rect 333716 122602 333744 124100
rect 344296 122602 344324 146270
rect 345018 133648 345074 133657
rect 345018 133583 345074 133592
rect 345032 125526 345060 133583
rect 345020 125520 345072 125526
rect 345020 125462 345072 125468
rect 345676 124846 345704 146406
rect 352012 146396 352064 146402
rect 352012 146338 352064 146344
rect 352024 143956 352052 146338
rect 361684 143956 361712 146406
rect 371332 146328 371384 146334
rect 371332 146270 371384 146276
rect 371344 143956 371372 146270
rect 350446 134328 350502 134337
rect 350446 134263 350502 134272
rect 350460 125526 350488 134263
rect 350448 125520 350500 125526
rect 350448 125462 350500 125468
rect 345664 124840 345716 124846
rect 371528 124794 371556 146406
rect 374644 146396 374696 146402
rect 374644 146338 374696 146344
rect 373264 146328 373316 146334
rect 373264 146270 373316 146276
rect 345664 124782 345716 124788
rect 371358 124766 371556 124794
rect 352024 122670 352052 124100
rect 361684 122670 361712 124100
rect 373276 122670 373304 146270
rect 373998 133648 374054 133657
rect 373998 133583 374054 133592
rect 374012 125594 374040 133583
rect 374000 125588 374052 125594
rect 374000 125530 374052 125536
rect 374656 122806 374684 146338
rect 389376 143970 389404 146406
rect 399024 146328 399076 146334
rect 399024 146270 399076 146276
rect 399036 143970 399064 146270
rect 389376 143942 389712 143970
rect 399036 143942 399372 143970
rect 379624 143262 380052 143290
rect 378046 134328 378102 134337
rect 378046 134263 378102 134272
rect 378060 125458 378088 134263
rect 378048 125452 378100 125458
rect 378048 125394 378100 125400
rect 374644 122800 374696 122806
rect 374644 122742 374696 122748
rect 379624 122670 379652 143262
rect 399496 124794 399524 146406
rect 400864 146328 400916 146334
rect 400864 146270 400916 146276
rect 399372 124766 399524 124794
rect 379716 124086 380052 124114
rect 389712 124086 390048 124114
rect 379716 122806 379744 124086
rect 379704 122800 379756 122806
rect 379704 122742 379756 122748
rect 352012 122664 352064 122670
rect 352012 122606 352064 122612
rect 361672 122664 361724 122670
rect 361672 122606 361724 122612
rect 373264 122664 373316 122670
rect 373264 122606 373316 122612
rect 379612 122664 379664 122670
rect 379612 122606 379664 122612
rect 390020 122602 390048 124086
rect 400876 122602 400904 146270
rect 408052 143956 408080 146474
rect 417700 146464 417752 146470
rect 417700 146406 417752 146412
rect 417712 143956 417740 146406
rect 428464 146396 428516 146402
rect 428464 146338 428516 146344
rect 427360 146328 427412 146334
rect 427360 146270 427412 146276
rect 427372 143956 427400 146270
rect 405646 134328 405702 134337
rect 405646 134263 405702 134272
rect 401598 133648 401654 133657
rect 401598 133583 401654 133592
rect 401612 125526 401640 133583
rect 405660 125594 405688 134263
rect 428476 132494 428504 146338
rect 428556 146328 428608 146334
rect 428556 146270 428608 146276
rect 427832 132466 428504 132494
rect 405648 125588 405700 125594
rect 405648 125530 405700 125536
rect 401600 125520 401652 125526
rect 401600 125462 401652 125468
rect 427832 124794 427860 132466
rect 427386 124766 427860 124794
rect 408052 122670 408080 124100
rect 417712 122670 417740 124100
rect 428568 122670 428596 146270
rect 428660 126274 428688 146474
rect 456064 146464 456116 146470
rect 456064 146406 456116 146412
rect 473360 146464 473412 146470
rect 473360 146406 473412 146412
rect 483480 146464 483532 146470
rect 483480 146406 483532 146412
rect 445668 146396 445720 146402
rect 445668 146338 445720 146344
rect 445680 143956 445708 146338
rect 455328 146328 455380 146334
rect 455328 146270 455380 146276
rect 455340 143956 455368 146270
rect 434824 143262 436034 143290
rect 434626 134328 434682 134337
rect 434626 134263 434682 134272
rect 429198 133648 429254 133657
rect 429198 133583 429254 133592
rect 428648 126268 428700 126274
rect 428648 126210 428700 126216
rect 429212 125458 429240 133583
rect 434640 125526 434668 134263
rect 434628 125520 434680 125526
rect 434628 125462 434680 125468
rect 429200 125452 429252 125458
rect 429200 125394 429252 125400
rect 434824 122670 434852 143262
rect 456076 132494 456104 146406
rect 464344 146396 464396 146402
rect 464344 146338 464396 146344
rect 456156 146328 456208 146334
rect 456156 146270 456208 146276
rect 455800 132466 456104 132494
rect 435732 126268 435784 126274
rect 435732 126210 435784 126216
rect 435744 124794 435772 126210
rect 455800 124794 455828 132466
rect 435744 124766 436034 124794
rect 455354 124766 455828 124794
rect 408040 122664 408092 122670
rect 408040 122606 408092 122612
rect 417700 122664 417752 122670
rect 417700 122606 417752 122612
rect 428556 122664 428608 122670
rect 428556 122606 428608 122612
rect 434812 122664 434864 122670
rect 434812 122606 434864 122612
rect 445680 122602 445708 124100
rect 456168 122602 456196 146270
rect 464356 143970 464384 146338
rect 464048 143942 464384 143970
rect 473372 143970 473400 146406
rect 483020 146328 483072 146334
rect 483020 146270 483072 146276
rect 483032 143970 483060 146270
rect 473372 143942 473708 143970
rect 483032 143942 483368 143970
rect 462226 134328 462282 134337
rect 462226 134263 462282 134272
rect 458178 133648 458234 133657
rect 458178 133583 458234 133592
rect 458192 125594 458220 133583
rect 458180 125588 458232 125594
rect 458180 125530 458232 125536
rect 462240 125458 462268 134263
rect 462228 125452 462280 125458
rect 462228 125394 462280 125400
rect 483492 124794 483520 146406
rect 483664 146396 483716 146402
rect 483664 146338 483716 146344
rect 483676 126954 483704 146338
rect 485044 146328 485096 146334
rect 485044 146270 485096 146276
rect 483664 126948 483716 126954
rect 483664 126890 483716 126896
rect 483368 124766 483520 124794
rect 463804 124086 464048 124114
rect 473708 124086 474044 124114
rect 463804 122670 463832 124086
rect 474016 122670 474044 124086
rect 485056 122670 485084 146270
rect 489826 134328 489882 134337
rect 489826 134263 489882 134272
rect 485778 133648 485834 133657
rect 485778 133583 485834 133592
rect 485792 125526 485820 133583
rect 489840 125594 489868 134263
rect 489828 125588 489880 125594
rect 489828 125530 489880 125536
rect 485780 125520 485832 125526
rect 485780 125462 485832 125468
rect 463792 122664 463844 122670
rect 463792 122606 463844 122612
rect 474004 122664 474056 122670
rect 474004 122606 474056 122612
rect 485044 122664 485096 122670
rect 485044 122606 485096 122612
rect 249708 122596 249760 122602
rect 249708 122538 249760 122544
rect 260196 122596 260248 122602
rect 260196 122538 260248 122544
rect 333704 122596 333756 122602
rect 333704 122538 333756 122544
rect 344284 122596 344336 122602
rect 344284 122538 344336 122544
rect 390008 122596 390060 122602
rect 390008 122538 390060 122544
rect 400864 122596 400916 122602
rect 400864 122538 400916 122544
rect 445668 122596 445720 122602
rect 445668 122538 445720 122544
rect 456156 122596 456208 122602
rect 456156 122538 456208 122544
rect 261484 118992 261536 118998
rect 261484 118934 261536 118940
rect 249708 118856 249760 118862
rect 249708 118798 249760 118804
rect 260104 118856 260156 118862
rect 260104 118798 260156 118804
rect 249720 116892 249748 118798
rect 259368 118788 259420 118794
rect 259368 118730 259420 118736
rect 259380 116892 259408 118730
rect 238864 116334 240074 116362
rect 238666 107264 238722 107273
rect 238666 107199 238722 107208
rect 238680 97918 238708 107199
rect 238668 97912 238720 97918
rect 238668 97854 238720 97860
rect 238864 95062 238892 116334
rect 260116 103514 260144 118798
rect 260196 118720 260248 118726
rect 260196 118662 260248 118668
rect 259840 103486 260144 103514
rect 239772 98252 239824 98258
rect 239772 98194 239824 98200
rect 239784 97730 239812 98194
rect 259840 97730 259868 103486
rect 239784 97702 240074 97730
rect 259394 97702 259868 97730
rect 238852 95056 238904 95062
rect 238852 94998 238904 95004
rect 249720 94994 249748 97036
rect 260208 94994 260236 118662
rect 249708 94988 249760 94994
rect 249708 94930 249760 94936
rect 260196 94988 260248 94994
rect 260196 94930 260248 94936
rect 260196 91248 260248 91254
rect 260196 91190 260248 91196
rect 249708 91180 249760 91186
rect 249708 91122 249760 91128
rect 249720 89964 249748 91122
rect 259368 91112 259420 91118
rect 259368 91054 259420 91060
rect 260104 91112 260156 91118
rect 260104 91054 260156 91060
rect 259380 89964 259408 91054
rect 238864 89270 240074 89298
rect 238668 88460 238720 88466
rect 238668 88402 238720 88408
rect 238680 80345 238708 88402
rect 238666 80336 238722 80345
rect 238666 80271 238722 80280
rect 238864 68882 238892 89270
rect 239772 72344 239824 72350
rect 239772 72286 239824 72292
rect 259736 72344 259788 72350
rect 259736 72286 259788 72292
rect 239784 70666 239812 72286
rect 259748 70666 259776 72286
rect 239784 70638 240074 70666
rect 259394 70638 259776 70666
rect 249720 68950 249748 70108
rect 260116 68950 260144 91054
rect 260208 72350 260236 91190
rect 260196 72344 260248 72350
rect 260196 72286 260248 72292
rect 261496 68950 261524 118934
rect 408040 118924 408092 118930
rect 408040 118866 408092 118872
rect 428648 118924 428700 118930
rect 428648 118866 428700 118872
rect 277676 118856 277728 118862
rect 277676 118798 277728 118804
rect 287520 118856 287572 118862
rect 287520 118798 287572 118804
rect 305368 118856 305420 118862
rect 305368 118798 305420 118804
rect 315488 118856 315540 118862
rect 315488 118798 315540 118804
rect 333704 118856 333756 118862
rect 333704 118798 333756 118804
rect 345664 118856 345716 118862
rect 345664 118798 345716 118804
rect 361672 118856 361724 118862
rect 361672 118798 361724 118804
rect 371516 118856 371568 118862
rect 371516 118798 371568 118804
rect 389364 118856 389416 118862
rect 389364 118798 389416 118804
rect 399484 118856 399536 118862
rect 399484 118798 399536 118804
rect 268016 118788 268068 118794
rect 268016 118730 268068 118736
rect 268028 116892 268056 118730
rect 277688 116892 277716 118798
rect 287336 118720 287388 118726
rect 287336 118662 287388 118668
rect 287348 116892 287376 118662
rect 266266 107264 266322 107273
rect 266266 107199 266322 107208
rect 262218 106584 262274 106593
rect 262218 106519 262274 106528
rect 262232 97986 262260 106519
rect 266280 97986 266308 107199
rect 262220 97980 262272 97986
rect 262220 97922 262272 97928
rect 266268 97980 266320 97986
rect 266268 97922 266320 97928
rect 287532 97730 287560 118798
rect 287704 118788 287756 118794
rect 287704 118730 287756 118736
rect 296352 118788 296404 118794
rect 296352 118730 296404 118736
rect 287716 98802 287744 118730
rect 289084 118720 289136 118726
rect 289084 118662 289136 118668
rect 287704 98796 287756 98802
rect 287704 98738 287756 98744
rect 287362 97702 287560 97730
rect 268028 95062 268056 97036
rect 277688 95062 277716 97036
rect 289096 95062 289124 118662
rect 296364 116906 296392 118730
rect 296056 116878 296392 116906
rect 305380 116906 305408 118798
rect 315028 118720 315080 118726
rect 315028 118662 315080 118668
rect 315040 116906 315068 118662
rect 305380 116878 305716 116906
rect 315040 116878 315376 116906
rect 293866 107264 293922 107273
rect 293866 107199 293922 107208
rect 289818 106584 289874 106593
rect 289818 106519 289874 106528
rect 289832 97918 289860 106519
rect 293880 97918 293908 107199
rect 295708 98796 295760 98802
rect 295708 98738 295760 98744
rect 289820 97912 289872 97918
rect 289820 97854 289872 97860
rect 293868 97912 293920 97918
rect 293868 97854 293920 97860
rect 295720 97730 295748 98738
rect 315500 97730 315528 118798
rect 316776 118788 316828 118794
rect 316776 118730 316828 118736
rect 316684 118720 316736 118726
rect 316684 118662 316736 118668
rect 295720 97702 296056 97730
rect 315376 97702 315528 97730
rect 305716 97022 306052 97050
rect 306024 95062 306052 97022
rect 316696 95062 316724 118662
rect 316788 98938 316816 118730
rect 333716 116892 333744 118798
rect 343364 118720 343416 118726
rect 343364 118662 343416 118668
rect 344284 118720 344336 118726
rect 344284 118662 344336 118668
rect 343376 116892 343404 118662
rect 323044 116334 324070 116362
rect 322846 107264 322902 107273
rect 322846 107199 322902 107208
rect 317418 106584 317474 106593
rect 317418 106519 317474 106528
rect 316776 98932 316828 98938
rect 316776 98874 316828 98880
rect 317432 97986 317460 106519
rect 322860 97986 322888 107199
rect 317420 97980 317472 97986
rect 317420 97922 317472 97928
rect 322848 97980 322900 97986
rect 322848 97922 322900 97928
rect 323044 95062 323072 116334
rect 323676 98932 323728 98938
rect 323676 98874 323728 98880
rect 323688 97730 323716 98874
rect 323688 97702 324070 97730
rect 343390 97714 343680 97730
rect 343390 97708 343692 97714
rect 343390 97702 343640 97708
rect 343640 97650 343692 97656
rect 268016 95056 268068 95062
rect 268016 94998 268068 95004
rect 277676 95056 277728 95062
rect 277676 94998 277728 95004
rect 289084 95056 289136 95062
rect 289084 94998 289136 95004
rect 306012 95056 306064 95062
rect 306012 94998 306064 95004
rect 316684 95056 316736 95062
rect 316684 94998 316736 95004
rect 323032 95056 323084 95062
rect 323032 94998 323084 95004
rect 333716 94994 333744 97036
rect 344296 94994 344324 118662
rect 345018 106584 345074 106593
rect 345018 106519 345074 106528
rect 345032 97918 345060 106519
rect 345020 97912 345072 97918
rect 345020 97854 345072 97860
rect 345676 97714 345704 118798
rect 352012 118788 352064 118794
rect 352012 118730 352064 118736
rect 352024 116892 352052 118730
rect 361684 116892 361712 118798
rect 371332 118720 371384 118726
rect 371332 118662 371384 118668
rect 371344 116892 371372 118662
rect 350446 107264 350502 107273
rect 350446 107199 350502 107208
rect 350460 97850 350488 107199
rect 350448 97844 350500 97850
rect 350448 97786 350500 97792
rect 371528 97730 371556 118798
rect 374644 118788 374696 118794
rect 374644 118730 374696 118736
rect 373264 118720 373316 118726
rect 373264 118662 373316 118668
rect 345664 97708 345716 97714
rect 371358 97702 371556 97730
rect 345664 97650 345716 97656
rect 352024 95062 352052 97036
rect 361684 95062 361712 97036
rect 373276 95062 373304 118662
rect 373998 106584 374054 106593
rect 373998 106519 374054 106528
rect 374012 97986 374040 106519
rect 374000 97980 374052 97986
rect 374000 97922 374052 97928
rect 374656 95198 374684 118730
rect 389376 116906 389404 118798
rect 399024 118720 399076 118726
rect 399024 118662 399076 118668
rect 399036 116906 399064 118662
rect 389376 116878 389712 116906
rect 399036 116878 399372 116906
rect 379624 116334 380052 116362
rect 378046 107264 378102 107273
rect 378046 107199 378102 107208
rect 378060 97918 378088 107199
rect 378048 97912 378100 97918
rect 378048 97854 378100 97860
rect 374644 95192 374696 95198
rect 374644 95134 374696 95140
rect 379624 95062 379652 116334
rect 399496 97730 399524 118798
rect 400864 118720 400916 118726
rect 400864 118662 400916 118668
rect 399372 97702 399524 97730
rect 379716 97022 380052 97050
rect 389712 97022 390048 97050
rect 379716 95198 379744 97022
rect 379704 95192 379756 95198
rect 379704 95134 379756 95140
rect 352012 95056 352064 95062
rect 352012 94998 352064 95004
rect 361672 95056 361724 95062
rect 361672 94998 361724 95004
rect 373264 95056 373316 95062
rect 373264 94998 373316 95004
rect 379612 95056 379664 95062
rect 379612 94998 379664 95004
rect 390020 94994 390048 97022
rect 400876 94994 400904 118662
rect 408052 116892 408080 118866
rect 417700 118856 417752 118862
rect 417700 118798 417752 118804
rect 417712 116892 417740 118798
rect 428464 118788 428516 118794
rect 428464 118730 428516 118736
rect 427360 118720 427412 118726
rect 427360 118662 427412 118668
rect 427372 116892 427400 118662
rect 405646 107264 405702 107273
rect 405646 107199 405702 107208
rect 401598 106584 401654 106593
rect 401598 106519 401654 106528
rect 401612 97850 401640 106519
rect 405660 97986 405688 107199
rect 428476 103514 428504 118730
rect 428556 118720 428608 118726
rect 428556 118662 428608 118668
rect 427832 103486 428504 103514
rect 405648 97980 405700 97986
rect 405648 97922 405700 97928
rect 401600 97844 401652 97850
rect 401600 97786 401652 97792
rect 427832 97730 427860 103486
rect 427386 97702 427860 97730
rect 408052 95062 408080 97036
rect 417712 95062 417740 97036
rect 428568 95062 428596 118662
rect 428660 98666 428688 118866
rect 456156 118856 456208 118862
rect 456156 118798 456208 118804
rect 473360 118856 473412 118862
rect 473360 118798 473412 118804
rect 483480 118856 483532 118862
rect 483480 118798 483532 118804
rect 445668 118788 445720 118794
rect 445668 118730 445720 118736
rect 445680 116892 445708 118730
rect 455328 118720 455380 118726
rect 455328 118662 455380 118668
rect 456064 118720 456116 118726
rect 456064 118662 456116 118668
rect 455340 116892 455368 118662
rect 434824 116334 436034 116362
rect 434626 107264 434682 107273
rect 434626 107199 434682 107208
rect 429198 106584 429254 106593
rect 429198 106519 429254 106528
rect 428648 98660 428700 98666
rect 428648 98602 428700 98608
rect 429212 97918 429240 106519
rect 429200 97912 429252 97918
rect 429200 97854 429252 97860
rect 434640 97850 434668 107199
rect 434628 97844 434680 97850
rect 434628 97786 434680 97792
rect 434824 95062 434852 116334
rect 455696 100292 455748 100298
rect 455696 100234 455748 100240
rect 435732 98660 435784 98666
rect 435732 98602 435784 98608
rect 435744 97730 435772 98602
rect 455708 97730 455736 100234
rect 435744 97702 436034 97730
rect 455354 97702 455736 97730
rect 408040 95056 408092 95062
rect 408040 94998 408092 95004
rect 417700 95056 417752 95062
rect 417700 94998 417752 95004
rect 428556 95056 428608 95062
rect 428556 94998 428608 95004
rect 434812 95056 434864 95062
rect 434812 94998 434864 95004
rect 445680 94994 445708 97036
rect 456076 94994 456104 118662
rect 456168 100298 456196 118798
rect 464344 118788 464396 118794
rect 464344 118730 464396 118736
rect 464356 116906 464384 118730
rect 464048 116878 464384 116906
rect 473372 116906 473400 118798
rect 483020 118720 483072 118726
rect 483020 118662 483072 118668
rect 483032 116906 483060 118662
rect 473372 116878 473708 116906
rect 483032 116878 483368 116906
rect 462226 107264 462282 107273
rect 462226 107199 462282 107208
rect 458178 106584 458234 106593
rect 458178 106519 458234 106528
rect 456156 100292 456208 100298
rect 456156 100234 456208 100240
rect 458192 97986 458220 106519
rect 458180 97980 458232 97986
rect 458180 97922 458232 97928
rect 462240 97918 462268 107199
rect 462228 97912 462280 97918
rect 462228 97854 462280 97860
rect 483492 97730 483520 118798
rect 483664 118788 483716 118794
rect 483664 118730 483716 118736
rect 483676 98666 483704 118730
rect 485044 118720 485096 118726
rect 485044 118662 485096 118668
rect 483664 98660 483716 98666
rect 483664 98602 483716 98608
rect 483368 97702 483520 97730
rect 463712 97022 464048 97050
rect 473708 97022 474044 97050
rect 463712 95062 463740 97022
rect 474016 95062 474044 97022
rect 485056 95062 485084 118662
rect 489826 107264 489882 107273
rect 489826 107199 489882 107208
rect 485778 106584 485834 106593
rect 485778 106519 485834 106528
rect 485792 97850 485820 106519
rect 489840 97986 489868 107199
rect 489828 97980 489880 97986
rect 489828 97922 489880 97928
rect 485780 97844 485832 97850
rect 485780 97786 485832 97792
rect 463700 95056 463752 95062
rect 463700 94998 463752 95004
rect 474004 95056 474056 95062
rect 474004 94998 474056 95004
rect 485044 95056 485096 95062
rect 485044 94998 485096 95004
rect 333704 94988 333756 94994
rect 333704 94930 333756 94936
rect 344284 94988 344336 94994
rect 344284 94930 344336 94936
rect 390008 94988 390060 94994
rect 390008 94930 390060 94936
rect 400864 94988 400916 94994
rect 400864 94930 400916 94936
rect 445668 94988 445720 94994
rect 445668 94930 445720 94936
rect 456064 94988 456116 94994
rect 456064 94930 456116 94936
rect 296352 91316 296404 91322
rect 296352 91258 296404 91264
rect 316776 91316 316828 91322
rect 316776 91258 316828 91264
rect 408040 91316 408092 91322
rect 408040 91258 408092 91264
rect 428648 91316 428700 91322
rect 428648 91258 428700 91264
rect 277676 91248 277728 91254
rect 277676 91190 277728 91196
rect 287520 91248 287572 91254
rect 287520 91190 287572 91196
rect 268016 91180 268068 91186
rect 268016 91122 268068 91128
rect 268028 89964 268056 91122
rect 277688 89964 277716 91190
rect 287336 91112 287388 91118
rect 287336 91054 287388 91060
rect 287348 89964 287376 91054
rect 262220 88392 262272 88398
rect 262220 88334 262272 88340
rect 262232 79665 262260 88334
rect 266266 80336 266322 80345
rect 266266 80271 266322 80280
rect 262218 79656 262274 79665
rect 262218 79591 262274 79600
rect 266280 71738 266308 80271
rect 266268 71732 266320 71738
rect 266268 71674 266320 71680
rect 287532 70666 287560 91190
rect 287704 91180 287756 91186
rect 287704 91122 287756 91128
rect 287716 72146 287744 91122
rect 289084 91112 289136 91118
rect 289084 91054 289136 91060
rect 287704 72140 287756 72146
rect 287704 72082 287756 72088
rect 287362 70638 287560 70666
rect 249708 68944 249760 68950
rect 249708 68886 249760 68892
rect 260104 68944 260156 68950
rect 260104 68886 260156 68892
rect 261484 68944 261536 68950
rect 261484 68886 261536 68892
rect 268028 68882 268056 70108
rect 277688 68882 277716 70108
rect 289096 68882 289124 91054
rect 296364 89978 296392 91258
rect 305368 91248 305420 91254
rect 305368 91190 305420 91196
rect 296056 89950 296392 89978
rect 305380 89978 305408 91190
rect 315488 91180 315540 91186
rect 315488 91122 315540 91128
rect 315028 91112 315080 91118
rect 315028 91054 315080 91060
rect 315040 89978 315068 91054
rect 305380 89950 305716 89978
rect 315040 89950 315376 89978
rect 289820 88460 289872 88466
rect 289820 88402 289872 88408
rect 293868 88460 293920 88466
rect 293868 88402 293920 88408
rect 289832 79665 289860 88402
rect 293880 80345 293908 88402
rect 293866 80336 293922 80345
rect 293866 80271 293922 80280
rect 289818 79656 289874 79665
rect 289818 79591 289874 79600
rect 295708 72140 295760 72146
rect 295708 72082 295760 72088
rect 295720 70666 295748 72082
rect 315500 70666 315528 91122
rect 316684 91112 316736 91118
rect 316684 91054 316736 91060
rect 295720 70638 296056 70666
rect 315376 70638 315528 70666
rect 305716 70094 306052 70122
rect 306024 68882 306052 70094
rect 316696 68882 316724 91054
rect 316788 72350 316816 91258
rect 345664 91248 345716 91254
rect 345664 91190 345716 91196
rect 361672 91248 361724 91254
rect 361672 91190 361724 91196
rect 371516 91248 371568 91254
rect 371516 91190 371568 91196
rect 389364 91248 389416 91254
rect 389364 91190 389416 91196
rect 399484 91248 399536 91254
rect 399484 91190 399536 91196
rect 333704 91180 333756 91186
rect 333704 91122 333756 91128
rect 333716 89964 333744 91122
rect 343364 91112 343416 91118
rect 343364 91054 343416 91060
rect 344284 91112 344336 91118
rect 344284 91054 344336 91060
rect 343376 89964 343404 91054
rect 323044 89270 324070 89298
rect 322848 88392 322900 88398
rect 322848 88334 322900 88340
rect 322860 80345 322888 88334
rect 322846 80336 322902 80345
rect 322846 80271 322902 80280
rect 317418 79656 317474 79665
rect 317418 79591 317474 79600
rect 316776 72344 316828 72350
rect 316776 72286 316828 72292
rect 317432 71738 317460 79591
rect 317420 71732 317472 71738
rect 317420 71674 317472 71680
rect 323044 68882 323072 89270
rect 323676 72344 323728 72350
rect 323676 72286 323728 72292
rect 323688 70666 323716 72286
rect 343548 71732 343600 71738
rect 343548 71674 343600 71680
rect 343560 70666 343588 71674
rect 323688 70638 324070 70666
rect 343390 70638 343588 70666
rect 238852 68876 238904 68882
rect 238852 68818 238904 68824
rect 268016 68876 268068 68882
rect 268016 68818 268068 68824
rect 277676 68876 277728 68882
rect 277676 68818 277728 68824
rect 289084 68876 289136 68882
rect 289084 68818 289136 68824
rect 306012 68876 306064 68882
rect 306012 68818 306064 68824
rect 316684 68876 316736 68882
rect 316684 68818 316736 68824
rect 323032 68876 323084 68882
rect 323032 68818 323084 68824
rect 333716 68814 333744 70108
rect 344296 68814 344324 91054
rect 345020 88460 345072 88466
rect 345020 88402 345072 88408
rect 345032 79665 345060 88402
rect 345018 79656 345074 79665
rect 345018 79591 345074 79600
rect 345676 71738 345704 91190
rect 352012 91180 352064 91186
rect 352012 91122 352064 91128
rect 352024 89964 352052 91122
rect 361684 89964 361712 91190
rect 371332 91112 371384 91118
rect 371332 91054 371384 91060
rect 371344 89964 371372 91054
rect 350448 88460 350500 88466
rect 350448 88402 350500 88408
rect 350460 80345 350488 88402
rect 350446 80336 350502 80345
rect 350446 80271 350502 80280
rect 345664 71732 345716 71738
rect 345664 71674 345716 71680
rect 371528 70666 371556 91190
rect 374644 91180 374696 91186
rect 374644 91122 374696 91128
rect 373264 91112 373316 91118
rect 373264 91054 373316 91060
rect 371358 70638 371556 70666
rect 352024 68882 352052 70108
rect 361684 68882 361712 70108
rect 373276 68882 373304 91054
rect 374000 88392 374052 88398
rect 374000 88334 374052 88340
rect 374012 79665 374040 88334
rect 373998 79656 374054 79665
rect 373998 79591 374054 79600
rect 374656 69018 374684 91122
rect 389376 89978 389404 91190
rect 399024 91112 399076 91118
rect 399024 91054 399076 91060
rect 399036 89978 399064 91054
rect 389376 89950 389712 89978
rect 399036 89950 399372 89978
rect 379624 89270 380052 89298
rect 378046 80336 378102 80345
rect 378046 80271 378102 80280
rect 378060 71738 378088 80271
rect 378048 71732 378100 71738
rect 378048 71674 378100 71680
rect 374644 69012 374696 69018
rect 374644 68954 374696 68960
rect 379624 68882 379652 89270
rect 399496 70666 399524 91190
rect 400864 91112 400916 91118
rect 400864 91054 400916 91060
rect 399372 70638 399524 70666
rect 379716 70094 380052 70122
rect 389712 70094 390048 70122
rect 379716 69018 379744 70094
rect 379704 69012 379756 69018
rect 379704 68954 379756 68960
rect 352012 68876 352064 68882
rect 352012 68818 352064 68824
rect 361672 68876 361724 68882
rect 361672 68818 361724 68824
rect 373264 68876 373316 68882
rect 373264 68818 373316 68824
rect 379612 68876 379664 68882
rect 379612 68818 379664 68824
rect 390020 68814 390048 70094
rect 400876 68814 400904 91054
rect 408052 89964 408080 91258
rect 417700 91248 417752 91254
rect 417700 91190 417752 91196
rect 417712 89964 417740 91190
rect 428464 91180 428516 91186
rect 428464 91122 428516 91128
rect 427360 91112 427412 91118
rect 427360 91054 427412 91060
rect 427372 89964 427400 91054
rect 401600 88460 401652 88466
rect 401600 88402 401652 88408
rect 401612 79665 401640 88402
rect 405648 88392 405700 88398
rect 405648 88334 405700 88340
rect 405660 80345 405688 88334
rect 405646 80336 405702 80345
rect 405646 80271 405702 80280
rect 401598 79656 401654 79665
rect 401598 79591 401654 79600
rect 428476 74534 428504 91122
rect 428556 91112 428608 91118
rect 428556 91054 428608 91060
rect 427832 74506 428504 74534
rect 427832 70666 427860 74506
rect 427386 70638 427860 70666
rect 408052 68882 408080 70108
rect 417712 68882 417740 70108
rect 428568 68882 428596 91054
rect 428660 72486 428688 91258
rect 456156 91248 456208 91254
rect 456156 91190 456208 91196
rect 473360 91248 473412 91254
rect 473360 91190 473412 91196
rect 483480 91248 483532 91254
rect 483480 91190 483532 91196
rect 445668 91180 445720 91186
rect 445668 91122 445720 91128
rect 445680 89964 445708 91122
rect 455328 91112 455380 91118
rect 455328 91054 455380 91060
rect 456064 91112 456116 91118
rect 456064 91054 456116 91060
rect 455340 89964 455368 91054
rect 434824 89270 436034 89298
rect 434628 88460 434680 88466
rect 434628 88402 434680 88408
rect 434640 80345 434668 88402
rect 434626 80336 434682 80345
rect 434626 80271 434682 80280
rect 429198 79656 429254 79665
rect 429198 79591 429254 79600
rect 428648 72480 428700 72486
rect 428648 72422 428700 72428
rect 429212 71738 429240 79591
rect 429200 71732 429252 71738
rect 429200 71674 429252 71680
rect 434824 68882 434852 89270
rect 435732 72480 435784 72486
rect 435732 72422 435784 72428
rect 435744 70666 435772 72422
rect 455696 72344 455748 72350
rect 455696 72286 455748 72292
rect 455708 70666 455736 72286
rect 435744 70638 436034 70666
rect 455354 70638 455736 70666
rect 408040 68876 408092 68882
rect 408040 68818 408092 68824
rect 417700 68876 417752 68882
rect 417700 68818 417752 68824
rect 428556 68876 428608 68882
rect 428556 68818 428608 68824
rect 434812 68876 434864 68882
rect 434812 68818 434864 68824
rect 445680 68814 445708 70108
rect 456076 68814 456104 91054
rect 456168 72350 456196 91190
rect 464344 91180 464396 91186
rect 464344 91122 464396 91128
rect 464356 89978 464384 91122
rect 464048 89950 464384 89978
rect 473372 89978 473400 91190
rect 483020 91112 483072 91118
rect 483020 91054 483072 91060
rect 483032 89978 483060 91054
rect 473372 89950 473708 89978
rect 483032 89950 483368 89978
rect 458180 88392 458232 88398
rect 458180 88334 458232 88340
rect 458192 79665 458220 88334
rect 462226 80336 462282 80345
rect 462226 80271 462282 80280
rect 458178 79656 458234 79665
rect 458178 79591 458234 79600
rect 456156 72344 456208 72350
rect 456156 72286 456208 72292
rect 462240 71670 462268 80271
rect 462228 71664 462280 71670
rect 462228 71606 462280 71612
rect 483492 70666 483520 91190
rect 483664 91180 483716 91186
rect 483664 91122 483716 91128
rect 483676 72282 483704 91122
rect 485044 91112 485096 91118
rect 485044 91054 485096 91060
rect 483664 72276 483716 72282
rect 483664 72218 483716 72224
rect 483368 70638 483520 70666
rect 463712 70094 464048 70122
rect 473708 70094 474044 70122
rect 463712 68882 463740 70094
rect 474016 68882 474044 70094
rect 485056 68882 485084 91054
rect 485780 88460 485832 88466
rect 485780 88402 485832 88408
rect 485792 79665 485820 88402
rect 489826 80336 489882 80345
rect 489826 80271 489882 80280
rect 485778 79656 485834 79665
rect 485778 79591 485834 79600
rect 489840 71738 489868 80271
rect 489828 71732 489880 71738
rect 489828 71674 489880 71680
rect 463700 68876 463752 68882
rect 463700 68818 463752 68824
rect 474004 68876 474056 68882
rect 474004 68818 474056 68824
rect 485044 68876 485096 68882
rect 485044 68818 485096 68824
rect 333704 68808 333756 68814
rect 333704 68750 333756 68756
rect 344284 68808 344336 68814
rect 344284 68750 344336 68756
rect 390008 68808 390060 68814
rect 390008 68750 390060 68756
rect 400864 68808 400916 68814
rect 400864 68750 400916 68756
rect 445668 68808 445720 68814
rect 445668 68750 445720 68756
rect 456064 68808 456116 68814
rect 456064 68750 456116 68756
rect 261484 65204 261536 65210
rect 261484 65146 261536 65152
rect 249708 65068 249760 65074
rect 249708 65010 249760 65016
rect 260104 65068 260156 65074
rect 260104 65010 260156 65016
rect 249720 62900 249748 65010
rect 259368 65000 259420 65006
rect 259368 64942 259420 64948
rect 259380 62900 259408 64942
rect 238864 62206 240074 62234
rect 238668 62144 238720 62150
rect 238668 62086 238720 62092
rect 238680 53281 238708 62086
rect 238666 53272 238722 53281
rect 238666 53207 238722 53216
rect 238864 41274 238892 62206
rect 260116 45554 260144 65010
rect 260196 64932 260248 64938
rect 260196 64874 260248 64880
rect 259840 45526 260144 45554
rect 239772 44940 239824 44946
rect 239772 44882 239824 44888
rect 239784 43738 239812 44882
rect 259840 43738 259868 45526
rect 239784 43710 240074 43738
rect 259394 43710 259868 43738
rect 238852 41268 238904 41274
rect 238852 41210 238904 41216
rect 249720 41206 249748 43044
rect 260208 41206 260236 64874
rect 249708 41200 249760 41206
rect 249708 41142 249760 41148
rect 260196 41200 260248 41206
rect 260196 41142 260248 41148
rect 234620 38072 234672 38078
rect 234620 38014 234672 38020
rect 212356 37528 212408 37534
rect 212356 37470 212408 37476
rect 232688 37528 232740 37534
rect 232688 37470 232740 37476
rect 148324 37460 148376 37466
rect 148324 37402 148376 37408
rect 165712 37460 165764 37466
rect 165712 37402 165764 37408
rect 175464 37460 175516 37466
rect 175464 37402 175516 37408
rect 193680 37460 193732 37466
rect 193680 37402 193732 37408
rect 203524 37460 203576 37466
rect 203524 37402 203576 37408
rect 81440 37392 81492 37398
rect 81440 37334 81492 37340
rect 91468 37392 91520 37398
rect 91468 37334 91520 37340
rect 109684 37392 109736 37398
rect 109684 37334 109736 37340
rect 126244 37392 126296 37398
rect 126244 37334 126296 37340
rect 137652 37392 137704 37398
rect 137652 37334 137704 37340
rect 81452 35986 81480 37334
rect 91100 37324 91152 37330
rect 91100 37266 91152 37272
rect 91112 35986 91140 37266
rect 81452 35958 81696 35986
rect 91112 35958 91356 35986
rect 71884 35278 72036 35306
rect 70308 34536 70360 34542
rect 70308 34478 70360 34484
rect 68284 27600 68336 27606
rect 68284 27542 68336 27548
rect 70320 26897 70348 34478
rect 70306 26888 70362 26897
rect 70306 26823 70362 26832
rect 65524 13796 65576 13802
rect 65524 13738 65576 13744
rect 64328 13660 64380 13666
rect 64328 13602 64380 13608
rect 71884 13530 71912 35278
rect 91480 16674 91508 37334
rect 93124 37324 93176 37330
rect 93124 37266 93176 37272
rect 91356 16646 91508 16674
rect 72036 16102 72096 16130
rect 81696 16102 82032 16130
rect 71872 13524 71924 13530
rect 71872 13466 71924 13472
rect 72068 13462 72096 16102
rect 82004 13802 82032 16102
rect 93136 13802 93164 37266
rect 93860 36032 93912 36038
rect 93860 35974 93912 35980
rect 93872 25673 93900 35974
rect 109696 35972 109724 37334
rect 119344 37324 119396 37330
rect 119344 37266 119396 37272
rect 120724 37324 120776 37330
rect 120724 37266 120776 37272
rect 119356 35972 119384 37266
rect 99484 35278 100050 35306
rect 97908 34604 97960 34610
rect 97908 34546 97960 34552
rect 97920 26353 97948 34546
rect 97906 26344 97962 26353
rect 97906 26279 97962 26288
rect 93858 25664 93914 25673
rect 93858 25599 93914 25608
rect 81992 13796 82044 13802
rect 81992 13738 82044 13744
rect 93124 13796 93176 13802
rect 93124 13738 93176 13744
rect 99484 13462 99512 35278
rect 100036 13530 100064 16116
rect 109696 13734 109724 16116
rect 119356 13802 119384 16116
rect 119344 13796 119396 13802
rect 119344 13738 119396 13744
rect 120736 13734 120764 37266
rect 121460 34536 121512 34542
rect 121460 34478 121512 34484
rect 121472 25673 121500 34478
rect 121458 25664 121514 25673
rect 121458 25599 121514 25608
rect 126256 13802 126284 37334
rect 137664 35972 137692 37334
rect 147312 37324 147364 37330
rect 147312 37266 147364 37272
rect 147324 35972 147352 37266
rect 127084 35278 128018 35306
rect 126888 34672 126940 34678
rect 126888 34614 126940 34620
rect 126900 26353 126928 34614
rect 126886 26344 126942 26353
rect 126886 26279 126942 26288
rect 126244 13796 126296 13802
rect 126244 13738 126296 13744
rect 109684 13728 109736 13734
rect 109684 13670 109736 13676
rect 120724 13728 120776 13734
rect 120724 13670 120776 13676
rect 100024 13524 100076 13530
rect 100024 13466 100076 13472
rect 127084 13462 127112 35278
rect 148336 16574 148364 37402
rect 156328 37392 156380 37398
rect 156328 37334 156380 37340
rect 148416 37324 148468 37330
rect 148416 37266 148468 37272
rect 147784 16546 148364 16574
rect 147784 16538 147812 16546
rect 147338 16510 147812 16538
rect 128004 13530 128032 16116
rect 137664 13734 137692 16116
rect 148428 13734 148456 37266
rect 156340 35986 156368 37334
rect 165724 35986 165752 37402
rect 175372 37324 175424 37330
rect 175372 37266 175424 37272
rect 175384 35986 175412 37266
rect 156032 35958 156368 35986
rect 165692 35958 165752 35986
rect 175352 35958 175412 35986
rect 149060 34604 149112 34610
rect 149060 34546 149112 34552
rect 149072 25673 149100 34546
rect 154488 34536 154540 34542
rect 154488 34478 154540 34484
rect 154500 26353 154528 34478
rect 154486 26344 154542 26353
rect 154486 26279 154542 26288
rect 149058 25664 149114 25673
rect 149058 25599 149114 25608
rect 175476 16674 175504 37402
rect 178684 37392 178736 37398
rect 178684 37334 178736 37340
rect 177304 37324 177356 37330
rect 177304 37266 177356 37272
rect 175352 16646 175504 16674
rect 156032 16102 156092 16130
rect 165692 16102 166028 16130
rect 137652 13728 137704 13734
rect 137652 13670 137704 13676
rect 148416 13728 148468 13734
rect 148416 13670 148468 13676
rect 156064 13530 156092 16102
rect 166000 13530 166028 16102
rect 177316 13530 177344 37266
rect 178040 34672 178092 34678
rect 178040 34614 178092 34620
rect 178052 25673 178080 34614
rect 178038 25664 178094 25673
rect 178038 25599 178094 25608
rect 178696 13802 178724 37334
rect 193692 35972 193720 37402
rect 203340 37324 203392 37330
rect 203340 37266 203392 37272
rect 203352 35972 203380 37266
rect 183664 35278 184046 35306
rect 182088 34604 182140 34610
rect 182088 34546 182140 34552
rect 182100 26353 182128 34546
rect 182086 26344 182142 26353
rect 182086 26279 182142 26288
rect 178684 13796 178736 13802
rect 178684 13738 178736 13744
rect 183664 13530 183692 35278
rect 203536 16674 203564 37402
rect 204904 37324 204956 37330
rect 204904 37266 204956 37272
rect 203366 16646 203564 16674
rect 184032 13802 184060 16116
rect 193692 13802 193720 16116
rect 204916 13802 204944 37266
rect 212368 35986 212396 37470
rect 221372 37460 221424 37466
rect 221372 37402 221424 37408
rect 212060 35958 212396 35986
rect 221384 35986 221412 37402
rect 232596 37392 232648 37398
rect 232596 37334 232648 37340
rect 231032 37324 231084 37330
rect 231032 37266 231084 37272
rect 232504 37324 232556 37330
rect 232504 37266 232556 37272
rect 231044 35986 231072 37266
rect 221384 35958 221720 35986
rect 231044 35958 231380 35986
rect 205640 34536 205692 34542
rect 205640 34478 205692 34484
rect 209688 34536 209740 34542
rect 209688 34478 209740 34484
rect 205652 25945 205680 34478
rect 209700 26353 209728 34478
rect 209686 26344 209742 26353
rect 209686 26279 209742 26288
rect 205638 25936 205694 25945
rect 205638 25871 205694 25880
rect 231676 16584 231728 16590
rect 231380 16532 231676 16538
rect 231380 16526 231728 16532
rect 231380 16510 231716 16526
rect 211724 16102 212060 16130
rect 221720 16102 222056 16130
rect 184020 13796 184072 13802
rect 184020 13738 184072 13744
rect 193680 13796 193732 13802
rect 193680 13738 193732 13744
rect 204904 13796 204956 13802
rect 204904 13738 204956 13744
rect 211724 13530 211752 16102
rect 222028 13530 222056 16102
rect 232516 13530 232544 37266
rect 232608 16590 232636 37334
rect 232700 18018 232728 37470
rect 260196 37460 260248 37466
rect 260196 37402 260248 37408
rect 249708 37392 249760 37398
rect 249708 37334 249760 37340
rect 249720 35972 249748 37334
rect 259368 37324 259420 37330
rect 259368 37266 259420 37272
rect 260104 37324 260156 37330
rect 260104 37266 260156 37272
rect 259380 35972 259408 37266
rect 238864 35278 240074 35306
rect 233240 34604 233292 34610
rect 233240 34546 233292 34552
rect 238668 34604 238720 34610
rect 238668 34546 238720 34552
rect 233252 25673 233280 34546
rect 238680 26353 238708 34546
rect 238666 26344 238722 26353
rect 238666 26279 238722 26288
rect 233238 25664 233294 25673
rect 233238 25599 233294 25608
rect 232688 18012 232740 18018
rect 232688 17954 232740 17960
rect 232596 16584 232648 16590
rect 232596 16526 232648 16532
rect 127992 13524 128044 13530
rect 127992 13466 128044 13472
rect 156052 13524 156104 13530
rect 156052 13466 156104 13472
rect 165988 13524 166040 13530
rect 165988 13466 166040 13472
rect 177304 13524 177356 13530
rect 177304 13466 177356 13472
rect 183652 13524 183704 13530
rect 183652 13466 183704 13472
rect 211712 13524 211764 13530
rect 211712 13466 211764 13472
rect 222016 13524 222068 13530
rect 222016 13466 222068 13472
rect 232504 13524 232556 13530
rect 232504 13466 232556 13472
rect 238864 13462 238892 35278
rect 259736 21480 259788 21486
rect 259736 21422 259788 21428
rect 239772 18012 239824 18018
rect 239772 17954 239824 17960
rect 239784 16674 239812 17954
rect 259748 16674 259776 21422
rect 239784 16646 240074 16674
rect 259394 16646 259776 16674
rect 249720 13530 249748 16116
rect 260116 13530 260144 37266
rect 260208 21486 260236 37402
rect 260196 21480 260248 21486
rect 260196 21422 260248 21428
rect 261496 13530 261524 65146
rect 408040 65136 408092 65142
rect 408040 65078 408092 65084
rect 428648 65136 428700 65142
rect 428648 65078 428700 65084
rect 277676 65068 277728 65074
rect 277676 65010 277728 65016
rect 287520 65068 287572 65074
rect 287520 65010 287572 65016
rect 305368 65068 305420 65074
rect 305368 65010 305420 65016
rect 315488 65068 315540 65074
rect 315488 65010 315540 65016
rect 333704 65068 333756 65074
rect 333704 65010 333756 65016
rect 345664 65068 345716 65074
rect 345664 65010 345716 65016
rect 361672 65068 361724 65074
rect 361672 65010 361724 65016
rect 371516 65068 371568 65074
rect 371516 65010 371568 65016
rect 389364 65068 389416 65074
rect 389364 65010 389416 65016
rect 399484 65068 399536 65074
rect 399484 65010 399536 65016
rect 268016 65000 268068 65006
rect 268016 64942 268068 64948
rect 268028 62900 268056 64942
rect 277688 62900 277716 65010
rect 287336 64932 287388 64938
rect 287336 64874 287388 64880
rect 287348 62900 287376 64874
rect 266266 53272 266322 53281
rect 266266 53207 266322 53216
rect 262218 52592 262274 52601
rect 262218 52527 262274 52536
rect 262232 44130 262260 52527
rect 266280 44130 266308 53207
rect 262220 44124 262272 44130
rect 262220 44066 262272 44072
rect 266268 44124 266320 44130
rect 266268 44066 266320 44072
rect 287532 43738 287560 65010
rect 287704 65000 287756 65006
rect 287704 64942 287756 64948
rect 296352 65000 296404 65006
rect 296352 64942 296404 64948
rect 287716 44334 287744 64942
rect 289084 64932 289136 64938
rect 289084 64874 289136 64880
rect 287704 44328 287756 44334
rect 287704 44270 287756 44276
rect 287362 43710 287560 43738
rect 268028 41274 268056 43044
rect 277688 41274 277716 43044
rect 289096 41274 289124 64874
rect 296364 62914 296392 64942
rect 296056 62886 296392 62914
rect 305380 62914 305408 65010
rect 315028 64932 315080 64938
rect 315028 64874 315080 64880
rect 315040 62914 315068 64874
rect 305380 62886 305716 62914
rect 315040 62886 315376 62914
rect 289820 62144 289872 62150
rect 289820 62086 289872 62092
rect 293868 62144 293920 62150
rect 293868 62086 293920 62092
rect 289832 52601 289860 62086
rect 293880 53281 293908 62086
rect 293866 53272 293922 53281
rect 293866 53207 293922 53216
rect 289818 52592 289874 52601
rect 289818 52527 289874 52536
rect 295708 44328 295760 44334
rect 295708 44270 295760 44276
rect 295720 43738 295748 44270
rect 315500 43738 315528 65010
rect 316776 65000 316828 65006
rect 316776 64942 316828 64948
rect 316684 64932 316736 64938
rect 316684 64874 316736 64880
rect 295720 43710 296056 43738
rect 315376 43710 315528 43738
rect 305716 43030 306052 43058
rect 306024 41274 306052 43030
rect 316696 41274 316724 64874
rect 316788 44334 316816 64942
rect 333716 62900 333744 65010
rect 343364 64932 343416 64938
rect 343364 64874 343416 64880
rect 344284 64932 344336 64938
rect 344284 64874 344336 64880
rect 343376 62900 343404 64874
rect 323044 62206 324070 62234
rect 322846 53272 322902 53281
rect 322846 53207 322902 53216
rect 317418 52592 317474 52601
rect 317418 52527 317474 52536
rect 316776 44328 316828 44334
rect 316776 44270 316828 44276
rect 317432 44130 317460 52527
rect 322860 44130 322888 53207
rect 317420 44124 317472 44130
rect 317420 44066 317472 44072
rect 322848 44124 322900 44130
rect 322848 44066 322900 44072
rect 323044 41274 323072 62206
rect 323676 44328 323728 44334
rect 323676 44270 323728 44276
rect 323688 43738 323716 44270
rect 343548 44056 343600 44062
rect 343548 43998 343600 44004
rect 343560 43738 343588 43998
rect 323688 43710 324070 43738
rect 343390 43710 343588 43738
rect 268016 41268 268068 41274
rect 268016 41210 268068 41216
rect 277676 41268 277728 41274
rect 277676 41210 277728 41216
rect 289084 41268 289136 41274
rect 289084 41210 289136 41216
rect 306012 41268 306064 41274
rect 306012 41210 306064 41216
rect 316684 41268 316736 41274
rect 316684 41210 316736 41216
rect 323032 41268 323084 41274
rect 323032 41210 323084 41216
rect 333716 41206 333744 43044
rect 344296 41206 344324 64874
rect 345020 62144 345072 62150
rect 345020 62086 345072 62092
rect 345032 52601 345060 62086
rect 345018 52592 345074 52601
rect 345018 52527 345074 52536
rect 345676 44062 345704 65010
rect 352012 65000 352064 65006
rect 352012 64942 352064 64948
rect 352024 62900 352052 64942
rect 361684 62900 361712 65010
rect 371332 64932 371384 64938
rect 371332 64874 371384 64880
rect 371344 62900 371372 64874
rect 350448 62212 350500 62218
rect 350448 62154 350500 62160
rect 350460 53281 350488 62154
rect 350446 53272 350502 53281
rect 350446 53207 350502 53216
rect 345664 44056 345716 44062
rect 345664 43998 345716 44004
rect 371528 43738 371556 65010
rect 374644 65000 374696 65006
rect 374644 64942 374696 64948
rect 373264 64932 373316 64938
rect 373264 64874 373316 64880
rect 371358 43710 371556 43738
rect 352024 41274 352052 43044
rect 361684 41274 361712 43044
rect 373276 41274 373304 64874
rect 373998 52592 374054 52601
rect 373998 52527 374054 52536
rect 374012 44130 374040 52527
rect 374000 44124 374052 44130
rect 374000 44066 374052 44072
rect 374656 41410 374684 64942
rect 389376 62914 389404 65010
rect 399024 64932 399076 64938
rect 399024 64874 399076 64880
rect 399036 62914 399064 64874
rect 389376 62886 389712 62914
rect 399036 62886 399372 62914
rect 379624 62206 380052 62234
rect 378048 62144 378100 62150
rect 378048 62086 378100 62092
rect 378060 53281 378088 62086
rect 378046 53272 378102 53281
rect 378046 53207 378102 53216
rect 374644 41404 374696 41410
rect 374644 41346 374696 41352
rect 379624 41274 379652 62206
rect 399496 43738 399524 65010
rect 400864 64932 400916 64938
rect 400864 64874 400916 64880
rect 399372 43710 399524 43738
rect 379716 43030 380052 43058
rect 389712 43030 390048 43058
rect 379716 41410 379744 43030
rect 379704 41404 379756 41410
rect 379704 41346 379756 41352
rect 352012 41268 352064 41274
rect 352012 41210 352064 41216
rect 361672 41268 361724 41274
rect 361672 41210 361724 41216
rect 373264 41268 373316 41274
rect 373264 41210 373316 41216
rect 379612 41268 379664 41274
rect 379612 41210 379664 41216
rect 390020 41206 390048 43030
rect 400876 41206 400904 64874
rect 408052 62900 408080 65078
rect 417700 65068 417752 65074
rect 417700 65010 417752 65016
rect 417712 62900 417740 65010
rect 428464 65000 428516 65006
rect 428464 64942 428516 64948
rect 427360 64932 427412 64938
rect 427360 64874 427412 64880
rect 427372 62900 427400 64874
rect 401600 62212 401652 62218
rect 401600 62154 401652 62160
rect 401612 52601 401640 62154
rect 405646 53272 405702 53281
rect 405646 53207 405702 53216
rect 401598 52592 401654 52601
rect 401598 52527 401654 52536
rect 405660 44130 405688 53207
rect 428476 45554 428504 64942
rect 428556 64932 428608 64938
rect 428556 64874 428608 64880
rect 427832 45526 428504 45554
rect 405648 44124 405700 44130
rect 405648 44066 405700 44072
rect 427832 43738 427860 45526
rect 427386 43710 427860 43738
rect 408052 41274 408080 43044
rect 417712 41274 417740 43044
rect 428568 41274 428596 64874
rect 428660 44878 428688 65078
rect 456156 65068 456208 65074
rect 456156 65010 456208 65016
rect 473544 65068 473596 65074
rect 473544 65010 473596 65016
rect 483480 65068 483532 65074
rect 483480 65010 483532 65016
rect 445668 65000 445720 65006
rect 445668 64942 445720 64948
rect 445680 62900 445708 64942
rect 455328 64932 455380 64938
rect 455328 64874 455380 64880
rect 456064 64932 456116 64938
rect 456064 64874 456116 64880
rect 455340 62900 455368 64874
rect 434824 62206 436034 62234
rect 429200 62144 429252 62150
rect 429200 62086 429252 62092
rect 434628 62144 434680 62150
rect 434628 62086 434680 62092
rect 429212 52601 429240 62086
rect 434640 53281 434668 62086
rect 434626 53272 434682 53281
rect 434626 53207 434682 53216
rect 429198 52592 429254 52601
rect 429198 52527 429254 52536
rect 428648 44872 428700 44878
rect 428648 44814 428700 44820
rect 434824 41274 434852 62206
rect 455696 50380 455748 50386
rect 455696 50322 455748 50328
rect 435732 44872 435784 44878
rect 435732 44814 435784 44820
rect 435744 43738 435772 44814
rect 455708 43738 455736 50322
rect 435744 43710 436034 43738
rect 455354 43710 455736 43738
rect 408040 41268 408092 41274
rect 408040 41210 408092 41216
rect 417700 41268 417752 41274
rect 417700 41210 417752 41216
rect 428556 41268 428608 41274
rect 428556 41210 428608 41216
rect 434812 41268 434864 41274
rect 434812 41210 434864 41216
rect 445680 41206 445708 43044
rect 456076 41206 456104 64874
rect 456168 50386 456196 65010
rect 464344 65000 464396 65006
rect 464344 64942 464396 64948
rect 464356 62914 464384 64942
rect 464048 62886 464384 62914
rect 473556 62914 473584 65010
rect 483204 64932 483256 64938
rect 483204 64874 483256 64880
rect 483216 62914 483244 64874
rect 473556 62886 473708 62914
rect 483216 62886 483368 62914
rect 462226 53272 462282 53281
rect 462226 53207 462282 53216
rect 458178 52592 458234 52601
rect 458178 52527 458234 52536
rect 456156 50380 456208 50386
rect 456156 50322 456208 50328
rect 458192 44130 458220 52527
rect 462240 44130 462268 53207
rect 458180 44124 458232 44130
rect 458180 44066 458232 44072
rect 462228 44124 462280 44130
rect 462228 44066 462280 44072
rect 483492 43738 483520 65010
rect 483664 65000 483716 65006
rect 483664 64942 483716 64948
rect 483676 44674 483704 64942
rect 485044 64932 485096 64938
rect 485044 64874 485096 64880
rect 483664 44668 483716 44674
rect 483664 44610 483716 44616
rect 483368 43710 483520 43738
rect 463712 43030 464048 43058
rect 473708 43030 474044 43058
rect 463712 41274 463740 43030
rect 474016 41274 474044 43030
rect 485056 41274 485084 64874
rect 485780 62144 485832 62150
rect 485780 62086 485832 62092
rect 489828 62144 489880 62150
rect 489828 62086 489880 62092
rect 485792 52601 485820 62086
rect 489840 53281 489868 62086
rect 489826 53272 489882 53281
rect 489826 53207 489882 53216
rect 485778 52592 485834 52601
rect 485778 52527 485834 52536
rect 463700 41268 463752 41274
rect 463700 41210 463752 41216
rect 474004 41268 474056 41274
rect 474004 41210 474056 41216
rect 485044 41268 485096 41274
rect 485044 41210 485096 41216
rect 333704 41200 333756 41206
rect 333704 41142 333756 41148
rect 344284 41200 344336 41206
rect 344284 41142 344336 41148
rect 390008 41200 390060 41206
rect 390008 41142 390060 41148
rect 400864 41200 400916 41206
rect 400864 41142 400916 41148
rect 445668 41200 445720 41206
rect 445668 41142 445720 41148
rect 456064 41200 456116 41206
rect 456064 41142 456116 41148
rect 408040 37528 408092 37534
rect 408040 37470 408092 37476
rect 428648 37528 428700 37534
rect 428648 37470 428700 37476
rect 277676 37460 277728 37466
rect 277676 37402 277728 37408
rect 287520 37460 287572 37466
rect 287520 37402 287572 37408
rect 305368 37460 305420 37466
rect 305368 37402 305420 37408
rect 345664 37460 345716 37466
rect 345664 37402 345716 37408
rect 361672 37460 361724 37466
rect 361672 37402 361724 37408
rect 371516 37460 371568 37466
rect 371516 37402 371568 37408
rect 389364 37460 389416 37466
rect 389364 37402 389416 37408
rect 399484 37460 399536 37466
rect 399484 37402 399536 37408
rect 268016 37392 268068 37398
rect 268016 37334 268068 37340
rect 268028 35972 268056 37334
rect 277688 35972 277716 37402
rect 287336 37324 287388 37330
rect 287336 37266 287388 37272
rect 287348 35972 287376 37266
rect 262220 34536 262272 34542
rect 262220 34478 262272 34484
rect 266268 34536 266320 34542
rect 266268 34478 266320 34484
rect 262232 25673 262260 34478
rect 266280 26353 266308 34478
rect 266266 26344 266322 26353
rect 266266 26279 266322 26288
rect 262218 25664 262274 25673
rect 262218 25599 262274 25608
rect 287532 16674 287560 37402
rect 287704 37392 287756 37398
rect 287704 37334 287756 37340
rect 296168 37392 296220 37398
rect 296168 37334 296220 37340
rect 287716 18290 287744 37334
rect 289084 37324 289136 37330
rect 289084 37266 289136 37272
rect 287704 18284 287756 18290
rect 287704 18226 287756 18232
rect 287362 16646 287560 16674
rect 249708 13524 249760 13530
rect 249708 13466 249760 13472
rect 260104 13524 260156 13530
rect 260104 13466 260156 13472
rect 261484 13524 261536 13530
rect 261484 13466 261536 13472
rect 268028 13462 268056 16116
rect 277688 13802 277716 16116
rect 289096 13802 289124 37266
rect 296180 35986 296208 37334
rect 296056 35958 296208 35986
rect 305380 35986 305408 37402
rect 316776 37392 316828 37398
rect 316776 37334 316828 37340
rect 322204 37392 322256 37398
rect 322204 37334 322256 37340
rect 333704 37392 333756 37398
rect 333704 37334 333756 37340
rect 315028 37324 315080 37330
rect 315028 37266 315080 37272
rect 316684 37324 316736 37330
rect 316684 37266 316736 37272
rect 315040 35986 315068 37266
rect 305380 35958 305716 35986
rect 315040 35958 315376 35986
rect 289820 34604 289872 34610
rect 289820 34546 289872 34552
rect 293868 34604 293920 34610
rect 293868 34546 293920 34552
rect 289832 25673 289860 34546
rect 293880 26353 293908 34546
rect 293866 26344 293922 26353
rect 293866 26279 293922 26288
rect 289818 25664 289874 25673
rect 289818 25599 289874 25608
rect 295708 18284 295760 18290
rect 295708 18226 295760 18232
rect 295720 16674 295748 18226
rect 295720 16646 296056 16674
rect 305716 16102 306052 16130
rect 315376 16102 315712 16130
rect 277676 13796 277728 13802
rect 277676 13738 277728 13744
rect 289084 13796 289136 13802
rect 289084 13738 289136 13744
rect 306024 13734 306052 16102
rect 315684 13802 315712 16102
rect 315672 13796 315724 13802
rect 315672 13738 315724 13744
rect 316696 13734 316724 37266
rect 316788 18154 316816 37334
rect 317420 34536 317472 34542
rect 317420 34478 317472 34484
rect 317432 25673 317460 34478
rect 317418 25664 317474 25673
rect 317418 25599 317474 25608
rect 316776 18148 316828 18154
rect 316776 18090 316828 18096
rect 322216 13802 322244 37334
rect 333716 35972 333744 37334
rect 343364 37324 343416 37330
rect 343364 37266 343416 37272
rect 344284 37324 344336 37330
rect 344284 37266 344336 37272
rect 343376 35972 343404 37266
rect 323044 35278 324070 35306
rect 322848 34536 322900 34542
rect 322848 34478 322900 34484
rect 322860 26353 322888 34478
rect 322846 26344 322902 26353
rect 322846 26279 322902 26288
rect 322204 13796 322256 13802
rect 322204 13738 322256 13744
rect 306012 13728 306064 13734
rect 306012 13670 306064 13676
rect 316684 13728 316736 13734
rect 316684 13670 316736 13676
rect 323044 13462 323072 35278
rect 323676 18148 323728 18154
rect 323676 18090 323728 18096
rect 323688 16674 323716 18090
rect 323688 16646 324070 16674
rect 343548 16584 343600 16590
rect 343390 16532 343548 16538
rect 343390 16526 343600 16532
rect 343390 16510 343588 16526
rect 333716 13734 333744 16116
rect 344296 13734 344324 37266
rect 345020 34604 345072 34610
rect 345020 34546 345072 34552
rect 345032 25673 345060 34546
rect 345018 25664 345074 25673
rect 345018 25599 345074 25608
rect 345676 16590 345704 37402
rect 352012 37392 352064 37398
rect 352012 37334 352064 37340
rect 352024 35972 352052 37334
rect 361684 35972 361712 37402
rect 371332 37324 371384 37330
rect 371332 37266 371384 37272
rect 371344 35972 371372 37266
rect 350448 34672 350500 34678
rect 350448 34614 350500 34620
rect 350460 26353 350488 34614
rect 350446 26344 350502 26353
rect 350446 26279 350502 26288
rect 371528 16674 371556 37402
rect 374644 37392 374696 37398
rect 374644 37334 374696 37340
rect 373264 37324 373316 37330
rect 373264 37266 373316 37272
rect 371358 16646 371556 16674
rect 345664 16584 345716 16590
rect 345664 16526 345716 16532
rect 333704 13728 333756 13734
rect 333704 13670 333756 13676
rect 344284 13728 344336 13734
rect 344284 13670 344336 13676
rect 352024 13462 352052 16116
rect 361684 13802 361712 16116
rect 373276 13802 373304 37266
rect 374000 34536 374052 34542
rect 374000 34478 374052 34484
rect 374012 25673 374040 34478
rect 373998 25664 374054 25673
rect 373998 25599 374054 25608
rect 374656 13802 374684 37334
rect 389376 35986 389404 37402
rect 399024 37324 399076 37330
rect 399024 37266 399076 37272
rect 399036 35986 399064 37266
rect 389376 35958 389712 35986
rect 399036 35958 399372 35986
rect 379624 35278 380052 35306
rect 378048 34604 378100 34610
rect 378048 34546 378100 34552
rect 378060 26353 378088 34546
rect 378046 26344 378102 26353
rect 378046 26279 378102 26288
rect 361672 13796 361724 13802
rect 361672 13738 361724 13744
rect 373264 13796 373316 13802
rect 373264 13738 373316 13744
rect 374644 13796 374696 13802
rect 374644 13738 374696 13744
rect 379624 13462 379652 35278
rect 399496 16674 399524 37402
rect 400864 37324 400916 37330
rect 400864 37266 400916 37272
rect 399372 16646 399524 16674
rect 379716 16102 380052 16130
rect 389712 16102 390048 16130
rect 379716 13802 379744 16102
rect 390020 13802 390048 16102
rect 400876 13802 400904 37266
rect 408052 35972 408080 37470
rect 417700 37460 417752 37466
rect 417700 37402 417752 37408
rect 417712 35972 417740 37402
rect 428464 37392 428516 37398
rect 428464 37334 428516 37340
rect 427360 37324 427412 37330
rect 427360 37266 427412 37272
rect 427372 35972 427400 37266
rect 401600 34672 401652 34678
rect 401600 34614 401652 34620
rect 401612 25673 401640 34614
rect 405648 34536 405700 34542
rect 405648 34478 405700 34484
rect 405660 26353 405688 34478
rect 405646 26344 405702 26353
rect 405646 26279 405702 26288
rect 401598 25664 401654 25673
rect 401598 25599 401654 25608
rect 428476 16574 428504 37334
rect 428556 37324 428608 37330
rect 428556 37266 428608 37272
rect 427832 16546 428504 16574
rect 427832 16538 427860 16546
rect 427386 16510 427860 16538
rect 379704 13796 379756 13802
rect 379704 13738 379756 13744
rect 390008 13796 390060 13802
rect 390008 13738 390060 13744
rect 400864 13796 400916 13802
rect 400864 13738 400916 13744
rect 408052 13462 408080 16116
rect 417712 13734 417740 16116
rect 428568 13734 428596 37266
rect 428660 18630 428688 37470
rect 456064 37460 456116 37466
rect 456064 37402 456116 37408
rect 473360 37460 473412 37466
rect 473360 37402 473412 37408
rect 483480 37460 483532 37466
rect 483480 37402 483532 37408
rect 445668 37392 445720 37398
rect 445668 37334 445720 37340
rect 445680 35972 445708 37334
rect 455328 37324 455380 37330
rect 455328 37266 455380 37272
rect 455340 35972 455368 37266
rect 434824 35278 436034 35306
rect 434628 34672 434680 34678
rect 434628 34614 434680 34620
rect 429200 34604 429252 34610
rect 429200 34546 429252 34552
rect 429212 25673 429240 34546
rect 434640 26353 434668 34614
rect 434626 26344 434682 26353
rect 434626 26279 434682 26288
rect 429198 25664 429254 25673
rect 429198 25599 429254 25608
rect 428648 18624 428700 18630
rect 428648 18566 428700 18572
rect 417700 13728 417752 13734
rect 417700 13670 417752 13676
rect 428556 13728 428608 13734
rect 428556 13670 428608 13676
rect 434824 13462 434852 35278
rect 456076 26234 456104 37402
rect 464344 37392 464396 37398
rect 464344 37334 464396 37340
rect 456156 37324 456208 37330
rect 456156 37266 456208 37272
rect 455800 26206 456104 26234
rect 435732 18624 435784 18630
rect 435732 18566 435784 18572
rect 435744 16674 435772 18566
rect 455800 16674 455828 26206
rect 435744 16646 436034 16674
rect 455354 16646 455828 16674
rect 445680 13734 445708 16116
rect 456168 13734 456196 37266
rect 464356 35986 464384 37334
rect 464048 35958 464384 35986
rect 473372 35986 473400 37402
rect 483020 37324 483072 37330
rect 483020 37266 483072 37272
rect 483032 35986 483060 37266
rect 473372 35958 473708 35986
rect 483032 35958 483368 35986
rect 462228 34604 462280 34610
rect 462228 34546 462280 34552
rect 458180 34536 458232 34542
rect 458180 34478 458232 34484
rect 458192 25673 458220 34478
rect 462240 26353 462268 34546
rect 462226 26344 462282 26353
rect 462226 26279 462282 26288
rect 458178 25664 458234 25673
rect 458178 25599 458234 25608
rect 483492 16674 483520 37402
rect 483664 37392 483716 37398
rect 483664 37334 483716 37340
rect 483676 18018 483704 37334
rect 485044 37324 485096 37330
rect 485044 37266 485096 37272
rect 483664 18012 483716 18018
rect 483664 17954 483716 17960
rect 483368 16646 483520 16674
rect 463712 16102 464048 16130
rect 473708 16102 474044 16130
rect 445668 13728 445720 13734
rect 445668 13670 445720 13676
rect 456156 13728 456208 13734
rect 456156 13670 456208 13676
rect 463712 13462 463740 16102
rect 474016 13802 474044 16102
rect 485056 13802 485084 37266
rect 485780 34672 485832 34678
rect 485780 34614 485832 34620
rect 485792 25673 485820 34614
rect 489828 34536 489880 34542
rect 489828 34478 489880 34484
rect 489840 26353 489868 34478
rect 489826 26344 489882 26353
rect 489826 26279 489882 26288
rect 485778 25664 485834 25673
rect 485778 25599 485834 25608
rect 474004 13796 474056 13802
rect 474004 13738 474056 13744
rect 485044 13796 485096 13802
rect 485044 13738 485096 13744
rect 490576 13598 490604 699654
rect 492036 686112 492088 686118
rect 492036 686054 492088 686060
rect 512736 686112 512788 686118
rect 512736 686054 512788 686060
rect 492048 683876 492076 686054
rect 501696 686044 501748 686050
rect 501696 685986 501748 685992
rect 501708 683876 501736 685986
rect 511448 685976 511500 685982
rect 511448 685918 511500 685924
rect 511356 685908 511408 685914
rect 511356 685850 511408 685856
rect 511368 683876 511396 685850
rect 491668 665304 491720 665310
rect 491668 665246 491720 665252
rect 491680 664714 491708 665246
rect 511460 664714 511488 685918
rect 512644 685908 512696 685914
rect 512644 685850 512696 685856
rect 491680 664686 492062 664714
rect 511382 664686 511488 664714
rect 501708 662386 501736 664020
rect 512656 662386 512684 685850
rect 512748 665310 512776 686054
rect 529664 685976 529716 685982
rect 529664 685918 529716 685924
rect 543004 685976 543056 685982
rect 543004 685918 543056 685924
rect 557540 685976 557592 685982
rect 557540 685918 557592 685924
rect 529676 683876 529704 685918
rect 539324 685908 539376 685914
rect 539324 685850 539376 685856
rect 540244 685908 540296 685914
rect 540244 685850 540296 685856
rect 539336 683876 539364 685850
rect 519004 683318 520030 683346
rect 518806 674248 518862 674257
rect 518806 674183 518862 674192
rect 513378 673568 513434 673577
rect 513378 673503 513434 673512
rect 512736 665304 512788 665310
rect 512736 665246 512788 665252
rect 513392 665174 513420 673503
rect 518820 665174 518848 674183
rect 513380 665168 513432 665174
rect 513380 665110 513432 665116
rect 518808 665168 518860 665174
rect 518808 665110 518860 665116
rect 519004 662386 519032 683318
rect 519636 665304 519688 665310
rect 519636 665246 519688 665252
rect 519648 664714 519676 665246
rect 519648 664686 520030 664714
rect 501696 662380 501748 662386
rect 501696 662322 501748 662328
rect 512644 662380 512696 662386
rect 512644 662322 512696 662328
rect 518992 662380 519044 662386
rect 518992 662322 519044 662328
rect 529676 662250 529704 664020
rect 539336 662318 539364 664020
rect 539324 662312 539376 662318
rect 539324 662254 539376 662260
rect 540256 662250 540284 685850
rect 542360 683188 542412 683194
rect 542360 683130 542412 683136
rect 541624 673872 541676 673878
rect 541624 673814 541676 673820
rect 529664 662244 529716 662250
rect 529664 662186 529716 662192
rect 540244 662244 540296 662250
rect 540244 662186 540296 662192
rect 492036 658504 492088 658510
rect 492036 658446 492088 658452
rect 512736 658504 512788 658510
rect 512736 658446 512788 658452
rect 492048 656948 492076 658446
rect 501696 658436 501748 658442
rect 501696 658378 501748 658384
rect 501708 656948 501736 658378
rect 511448 658368 511500 658374
rect 511448 658310 511500 658316
rect 511356 658300 511408 658306
rect 511356 658242 511408 658248
rect 511368 656948 511396 658242
rect 491668 639396 491720 639402
rect 491668 639338 491720 639344
rect 491680 637786 491708 639338
rect 511460 637786 511488 658310
rect 512644 658300 512696 658306
rect 512644 658242 512696 658248
rect 491680 637758 492062 637786
rect 511382 637758 511488 637786
rect 501708 634642 501736 637092
rect 512656 634642 512684 658242
rect 512748 639130 512776 658446
rect 529664 658368 529716 658374
rect 529664 658310 529716 658316
rect 529676 656948 529704 658310
rect 539324 658300 539376 658306
rect 539324 658242 539376 658248
rect 540244 658300 540296 658306
rect 540244 658242 540296 658248
rect 539336 656948 539364 658242
rect 519004 656254 520030 656282
rect 513380 655716 513432 655722
rect 513380 655658 513432 655664
rect 513392 646649 513420 655658
rect 518808 655648 518860 655654
rect 518808 655590 518860 655596
rect 518820 647329 518848 655590
rect 518806 647320 518862 647329
rect 518806 647255 518862 647264
rect 513378 646640 513434 646649
rect 513378 646575 513434 646584
rect 512736 639124 512788 639130
rect 512736 639066 512788 639072
rect 519004 634642 519032 656254
rect 519636 639124 519688 639130
rect 519636 639066 519688 639072
rect 519648 637786 519676 639066
rect 519648 637758 520030 637786
rect 501696 634636 501748 634642
rect 501696 634578 501748 634584
rect 512644 634636 512696 634642
rect 512644 634578 512696 634584
rect 518992 634636 519044 634642
rect 518992 634578 519044 634584
rect 529676 634574 529704 637092
rect 539336 634778 539364 637092
rect 539324 634772 539376 634778
rect 539324 634714 539376 634720
rect 540256 634574 540284 658242
rect 529664 634568 529716 634574
rect 529664 634510 529716 634516
rect 540244 634568 540296 634574
rect 540244 634510 540296 634516
rect 492036 632324 492088 632330
rect 492036 632266 492088 632272
rect 512736 632324 512788 632330
rect 512736 632266 512788 632272
rect 492048 629884 492076 632266
rect 501696 632256 501748 632262
rect 501696 632198 501748 632204
rect 501708 629884 501736 632198
rect 511448 632188 511500 632194
rect 511448 632130 511500 632136
rect 511356 632120 511408 632126
rect 511356 632062 511408 632068
rect 511368 629884 511396 632062
rect 491668 611788 491720 611794
rect 491668 611730 491720 611736
rect 491680 610722 491708 611730
rect 511460 610722 511488 632130
rect 512644 632120 512696 632126
rect 512644 632062 512696 632068
rect 491680 610694 492062 610722
rect 511382 610694 511488 610722
rect 501708 608462 501736 610028
rect 512656 608462 512684 632062
rect 512748 611794 512776 632266
rect 529664 632188 529716 632194
rect 529664 632130 529716 632136
rect 529676 629884 529704 632130
rect 539324 632120 539376 632126
rect 539324 632062 539376 632068
rect 540244 632120 540296 632126
rect 540244 632062 540296 632068
rect 539336 629884 539364 632062
rect 519004 629326 520030 629354
rect 518806 620256 518862 620265
rect 518806 620191 518862 620200
rect 513378 619576 513434 619585
rect 513378 619511 513434 619520
rect 512736 611788 512788 611794
rect 512736 611730 512788 611736
rect 513392 611250 513420 619511
rect 518820 611250 518848 620191
rect 513380 611244 513432 611250
rect 513380 611186 513432 611192
rect 518808 611244 518860 611250
rect 518808 611186 518860 611192
rect 519004 608462 519032 629326
rect 519636 611788 519688 611794
rect 519636 611730 519688 611736
rect 519648 610722 519676 611730
rect 519648 610694 520030 610722
rect 501696 608456 501748 608462
rect 501696 608398 501748 608404
rect 512644 608456 512696 608462
rect 512644 608398 512696 608404
rect 518992 608456 519044 608462
rect 518992 608398 519044 608404
rect 529676 608394 529704 610028
rect 539336 608598 539364 610028
rect 539324 608592 539376 608598
rect 539324 608534 539376 608540
rect 540256 608394 540284 632062
rect 529664 608388 529716 608394
rect 529664 608330 529716 608336
rect 540244 608388 540296 608394
rect 540244 608330 540296 608336
rect 492036 604716 492088 604722
rect 492036 604658 492088 604664
rect 512736 604716 512788 604722
rect 512736 604658 512788 604664
rect 492048 602956 492076 604658
rect 501696 604648 501748 604654
rect 501696 604590 501748 604596
rect 501708 602956 501736 604590
rect 511448 604580 511500 604586
rect 511448 604522 511500 604528
rect 511356 604512 511408 604518
rect 511356 604454 511408 604460
rect 511368 602956 511396 604454
rect 491668 584180 491720 584186
rect 491668 584122 491720 584128
rect 491680 583794 491708 584122
rect 511460 583794 511488 604522
rect 512644 604512 512696 604518
rect 512644 604454 512696 604460
rect 491680 583766 492062 583794
rect 511382 583766 511488 583794
rect 501708 580854 501736 583100
rect 512656 580854 512684 604454
rect 512748 584322 512776 604658
rect 529664 604580 529716 604586
rect 529664 604522 529716 604528
rect 529676 602956 529704 604522
rect 539324 604512 539376 604518
rect 539324 604454 539376 604460
rect 540244 604512 540296 604518
rect 540244 604454 540296 604460
rect 539336 602956 539364 604454
rect 519004 602262 520030 602290
rect 518806 593328 518862 593337
rect 518806 593263 518862 593272
rect 513378 592648 513434 592657
rect 513378 592583 513434 592592
rect 512736 584316 512788 584322
rect 512736 584258 512788 584264
rect 513392 583574 513420 592583
rect 518820 583642 518848 593263
rect 518808 583636 518860 583642
rect 518808 583578 518860 583584
rect 513380 583568 513432 583574
rect 513380 583510 513432 583516
rect 519004 580854 519032 602262
rect 519636 584316 519688 584322
rect 519636 584258 519688 584264
rect 519648 583794 519676 584258
rect 519648 583766 520030 583794
rect 539508 583568 539560 583574
rect 539350 583516 539508 583522
rect 539350 583510 539560 583516
rect 539350 583494 539548 583510
rect 501696 580848 501748 580854
rect 501696 580790 501748 580796
rect 512644 580848 512696 580854
rect 512644 580790 512696 580796
rect 518992 580848 519044 580854
rect 518992 580790 519044 580796
rect 529676 580786 529704 583100
rect 540256 580786 540284 604454
rect 529664 580780 529716 580786
rect 529664 580722 529716 580728
rect 540244 580780 540296 580786
rect 540244 580722 540296 580728
rect 492036 578468 492088 578474
rect 492036 578410 492088 578416
rect 512736 578468 512788 578474
rect 512736 578410 512788 578416
rect 492048 575892 492076 578410
rect 501696 578400 501748 578406
rect 501696 578342 501748 578348
rect 501708 575892 501736 578342
rect 511448 578332 511500 578338
rect 511448 578274 511500 578280
rect 511356 578264 511408 578270
rect 511356 578206 511408 578212
rect 511368 575892 511396 578206
rect 491668 558204 491720 558210
rect 491668 558146 491720 558152
rect 491680 556730 491708 558146
rect 511460 556730 511488 578274
rect 512644 578264 512696 578270
rect 512644 578206 512696 578212
rect 491680 556702 492062 556730
rect 511382 556702 511488 556730
rect 501708 554606 501736 556036
rect 512656 554606 512684 578206
rect 512748 557666 512776 578410
rect 529664 578332 529716 578338
rect 529664 578274 529716 578280
rect 529676 575892 529704 578274
rect 539324 578264 539376 578270
rect 539324 578206 539376 578212
rect 540244 578264 540296 578270
rect 540244 578206 540296 578212
rect 539336 575892 539364 578206
rect 519004 575334 520030 575362
rect 518806 566264 518862 566273
rect 518806 566199 518862 566208
rect 513378 565584 513434 565593
rect 513378 565519 513434 565528
rect 512736 557660 512788 557666
rect 512736 557602 512788 557608
rect 513392 557394 513420 565519
rect 518820 557462 518848 566199
rect 518808 557456 518860 557462
rect 518808 557398 518860 557404
rect 513380 557388 513432 557394
rect 513380 557330 513432 557336
rect 519004 554606 519032 575334
rect 519636 557660 519688 557666
rect 519636 557602 519688 557608
rect 519648 556730 519676 557602
rect 519648 556702 520030 556730
rect 501696 554600 501748 554606
rect 501696 554542 501748 554548
rect 512644 554600 512696 554606
rect 512644 554542 512696 554548
rect 518992 554600 519044 554606
rect 518992 554542 519044 554548
rect 529676 554538 529704 556036
rect 539336 554742 539364 556036
rect 539324 554736 539376 554742
rect 539324 554678 539376 554684
rect 540256 554538 540284 578206
rect 529664 554532 529716 554538
rect 529664 554474 529716 554480
rect 540244 554532 540296 554538
rect 540244 554474 540296 554480
rect 492036 550860 492088 550866
rect 492036 550802 492088 550808
rect 512736 550860 512788 550866
rect 512736 550802 512788 550808
rect 492048 548964 492076 550802
rect 501696 550792 501748 550798
rect 501696 550734 501748 550740
rect 501708 548964 501736 550734
rect 511448 550724 511500 550730
rect 511448 550666 511500 550672
rect 511356 550656 511408 550662
rect 511356 550598 511408 550604
rect 511368 548964 511396 550598
rect 491668 530188 491720 530194
rect 491668 530130 491720 530136
rect 491680 529666 491708 530130
rect 511460 529666 511488 550666
rect 512644 550656 512696 550662
rect 512644 550598 512696 550604
rect 491680 529638 492062 529666
rect 511382 529638 511488 529666
rect 501708 526998 501736 529108
rect 512656 526998 512684 550598
rect 512748 530262 512776 550802
rect 529664 550724 529716 550730
rect 529664 550666 529716 550672
rect 529676 548964 529704 550666
rect 539324 550656 539376 550662
rect 539324 550598 539376 550604
rect 540244 550656 540296 550662
rect 540244 550598 540296 550604
rect 539336 548964 539364 550598
rect 519004 548270 520030 548298
rect 518806 539336 518862 539345
rect 518806 539271 518862 539280
rect 513378 538656 513434 538665
rect 513378 538591 513434 538600
rect 512736 530256 512788 530262
rect 512736 530198 512788 530204
rect 513392 529786 513420 538591
rect 518820 529854 518848 539271
rect 518808 529848 518860 529854
rect 518808 529790 518860 529796
rect 513380 529780 513432 529786
rect 513380 529722 513432 529728
rect 519004 526998 519032 548270
rect 519636 530256 519688 530262
rect 519636 530198 519688 530204
rect 519648 529666 519676 530198
rect 519648 529638 520030 529666
rect 501696 526992 501748 526998
rect 501696 526934 501748 526940
rect 512644 526992 512696 526998
rect 512644 526934 512696 526940
rect 518992 526992 519044 526998
rect 518992 526934 519044 526940
rect 529676 526930 529704 529108
rect 539336 527134 539364 529108
rect 539324 527128 539376 527134
rect 539324 527070 539376 527076
rect 540256 526930 540284 550598
rect 529664 526924 529716 526930
rect 529664 526866 529716 526872
rect 540244 526924 540296 526930
rect 540244 526866 540296 526872
rect 492036 523252 492088 523258
rect 492036 523194 492088 523200
rect 512736 523252 512788 523258
rect 512736 523194 512788 523200
rect 492048 521900 492076 523194
rect 501696 523184 501748 523190
rect 501696 523126 501748 523132
rect 501708 521900 501736 523126
rect 511448 523116 511500 523122
rect 511448 523058 511500 523064
rect 511356 523048 511408 523054
rect 511356 522990 511408 522996
rect 511368 521900 511396 522990
rect 491668 504348 491720 504354
rect 491668 504290 491720 504296
rect 491680 502738 491708 504290
rect 511460 502738 511488 523058
rect 512644 523048 512696 523054
rect 512644 522990 512696 522996
rect 491680 502710 492062 502738
rect 511382 502710 511488 502738
rect 501708 500818 501736 502044
rect 512656 500818 512684 522990
rect 512748 504354 512776 523194
rect 529664 523116 529716 523122
rect 529664 523058 529716 523064
rect 529676 521900 529704 523058
rect 539324 523048 539376 523054
rect 539324 522990 539376 522996
rect 540244 523048 540296 523054
rect 540244 522990 540296 522996
rect 539336 521900 539364 522990
rect 519004 521206 520030 521234
rect 518808 520328 518860 520334
rect 518808 520270 518860 520276
rect 518820 512281 518848 520270
rect 518806 512272 518862 512281
rect 518806 512207 518862 512216
rect 513378 511592 513434 511601
rect 513378 511527 513434 511536
rect 512736 504348 512788 504354
rect 512736 504290 512788 504296
rect 513392 503606 513420 511527
rect 513380 503600 513432 503606
rect 513380 503542 513432 503548
rect 519004 500818 519032 521206
rect 519636 504348 519688 504354
rect 519636 504290 519688 504296
rect 519648 502738 519676 504290
rect 519648 502710 520030 502738
rect 501696 500812 501748 500818
rect 501696 500754 501748 500760
rect 512644 500812 512696 500818
rect 512644 500754 512696 500760
rect 518992 500812 519044 500818
rect 518992 500754 519044 500760
rect 529676 500750 529704 502044
rect 539336 500954 539364 502044
rect 539324 500948 539376 500954
rect 539324 500890 539376 500896
rect 540256 500750 540284 522990
rect 540886 511048 540942 511057
rect 540886 510983 540942 510992
rect 540900 509250 540928 510983
rect 540888 509244 540940 509250
rect 540888 509186 540940 509192
rect 529664 500744 529716 500750
rect 529664 500686 529716 500692
rect 540244 500744 540296 500750
rect 540244 500686 540296 500692
rect 492036 497072 492088 497078
rect 492036 497014 492088 497020
rect 512736 497072 512788 497078
rect 512736 497014 512788 497020
rect 492048 494972 492076 497014
rect 501696 497004 501748 497010
rect 501696 496946 501748 496952
rect 501708 494972 501736 496946
rect 511448 496936 511500 496942
rect 511448 496878 511500 496884
rect 511356 496868 511408 496874
rect 511356 496810 511408 496816
rect 511368 494972 511396 496810
rect 491668 476332 491720 476338
rect 491668 476274 491720 476280
rect 491680 475674 491708 476274
rect 511460 475674 511488 496878
rect 512644 496868 512696 496874
rect 512644 496810 512696 496816
rect 491680 475646 492062 475674
rect 511382 475646 511488 475674
rect 501708 473210 501736 475116
rect 512656 473210 512684 496810
rect 512748 477018 512776 497014
rect 529664 496936 529716 496942
rect 529664 496878 529716 496884
rect 529676 494972 529704 496878
rect 539324 496868 539376 496874
rect 539324 496810 539376 496816
rect 540244 496868 540296 496874
rect 540244 496810 540296 496816
rect 539336 494972 539364 496810
rect 519004 494278 520030 494306
rect 518806 485344 518862 485353
rect 518806 485279 518862 485288
rect 513378 484664 513434 484673
rect 513378 484599 513434 484608
rect 512736 477012 512788 477018
rect 512736 476954 512788 476960
rect 513392 475930 513420 484599
rect 518820 475998 518848 485279
rect 518808 475992 518860 475998
rect 518808 475934 518860 475940
rect 513380 475924 513432 475930
rect 513380 475866 513432 475872
rect 519004 473210 519032 494278
rect 519636 477012 519688 477018
rect 519636 476954 519688 476960
rect 519648 475674 519676 476954
rect 539508 475924 539560 475930
rect 539508 475866 539560 475872
rect 539520 475674 539548 475866
rect 519648 475646 520030 475674
rect 539350 475646 539548 475674
rect 501696 473204 501748 473210
rect 501696 473146 501748 473152
rect 512644 473204 512696 473210
rect 512644 473146 512696 473152
rect 518992 473204 519044 473210
rect 518992 473146 519044 473152
rect 529676 473142 529704 475116
rect 540256 473142 540284 496810
rect 529664 473136 529716 473142
rect 529664 473078 529716 473084
rect 540244 473136 540296 473142
rect 540244 473078 540296 473084
rect 501696 469396 501748 469402
rect 501696 469338 501748 469344
rect 511448 469396 511500 469402
rect 511448 469338 511500 469344
rect 529664 469396 529716 469402
rect 529664 469338 529716 469344
rect 492036 469328 492088 469334
rect 492036 469270 492088 469276
rect 492048 467908 492076 469270
rect 501708 467908 501736 469338
rect 511356 469260 511408 469266
rect 511356 469202 511408 469208
rect 511368 467908 511396 469202
rect 491668 450356 491720 450362
rect 491668 450298 491720 450304
rect 491680 448746 491708 450298
rect 511460 448746 511488 469338
rect 512736 469328 512788 469334
rect 512736 469270 512788 469276
rect 512644 469260 512696 469266
rect 512644 469202 512696 469208
rect 491680 448718 492062 448746
rect 511382 448718 511488 448746
rect 501708 445602 501736 448052
rect 512656 445602 512684 469202
rect 512748 450498 512776 469270
rect 529676 467908 529704 469338
rect 539324 469260 539376 469266
rect 539324 469202 539376 469208
rect 540244 469260 540296 469266
rect 540244 469202 540296 469208
rect 539336 467908 539364 469202
rect 519004 467214 520030 467242
rect 513380 466608 513432 466614
rect 513380 466550 513432 466556
rect 513392 457609 513420 466550
rect 518808 466540 518860 466546
rect 518808 466482 518860 466488
rect 518820 458289 518848 466482
rect 518806 458280 518862 458289
rect 518806 458215 518862 458224
rect 513378 457600 513434 457609
rect 513378 457535 513434 457544
rect 512736 450492 512788 450498
rect 512736 450434 512788 450440
rect 519004 445602 519032 467214
rect 519636 450492 519688 450498
rect 519636 450434 519688 450440
rect 519648 448746 519676 450434
rect 519648 448718 520030 448746
rect 539508 448520 539560 448526
rect 539350 448468 539508 448474
rect 539350 448462 539560 448468
rect 539350 448446 539548 448462
rect 501696 445596 501748 445602
rect 501696 445538 501748 445544
rect 512644 445596 512696 445602
rect 512644 445538 512696 445544
rect 518992 445596 519044 445602
rect 518992 445538 519044 445544
rect 529676 445534 529704 448052
rect 540256 445534 540284 469202
rect 529664 445528 529716 445534
rect 529664 445470 529716 445476
rect 540244 445528 540296 445534
rect 540244 445470 540296 445476
rect 492036 443216 492088 443222
rect 492036 443158 492088 443164
rect 512736 443216 512788 443222
rect 512736 443158 512788 443164
rect 492048 440980 492076 443158
rect 501696 443148 501748 443154
rect 501696 443090 501748 443096
rect 501708 440980 501736 443090
rect 511448 443080 511500 443086
rect 511448 443022 511500 443028
rect 511356 443012 511408 443018
rect 511356 442954 511408 442960
rect 511368 440980 511396 442954
rect 491668 423088 491720 423094
rect 491668 423030 491720 423036
rect 491680 421682 491708 423030
rect 511460 421682 511488 443022
rect 512644 443012 512696 443018
rect 512644 442954 512696 442960
rect 491680 421654 492062 421682
rect 511382 421654 511488 421682
rect 501708 419354 501736 421124
rect 512656 419354 512684 442954
rect 512748 423026 512776 443158
rect 529664 443080 529716 443086
rect 529664 443022 529716 443028
rect 529676 440980 529704 443022
rect 539324 443012 539376 443018
rect 539324 442954 539376 442960
rect 540244 443012 540296 443018
rect 540244 442954 540296 442960
rect 539336 440980 539364 442954
rect 519004 440286 520030 440314
rect 518806 431352 518862 431361
rect 518806 431287 518862 431296
rect 513378 430672 513434 430681
rect 513378 430607 513434 430616
rect 512736 423020 512788 423026
rect 512736 422962 512788 422968
rect 513392 422278 513420 430607
rect 518820 422278 518848 431287
rect 513380 422272 513432 422278
rect 513380 422214 513432 422220
rect 518808 422272 518860 422278
rect 518808 422214 518860 422220
rect 519004 419354 519032 440286
rect 519636 423020 519688 423026
rect 519636 422962 519688 422968
rect 519648 421682 519676 422962
rect 539508 421728 539560 421734
rect 519648 421654 520030 421682
rect 539350 421676 539508 421682
rect 539350 421670 539560 421676
rect 539350 421654 539548 421670
rect 501696 419348 501748 419354
rect 501696 419290 501748 419296
rect 512644 419348 512696 419354
rect 512644 419290 512696 419296
rect 518992 419348 519044 419354
rect 518992 419290 519044 419296
rect 529676 419286 529704 421124
rect 540256 419286 540284 442954
rect 529664 419280 529716 419286
rect 529664 419222 529716 419228
rect 540244 419280 540296 419286
rect 540244 419222 540296 419228
rect 492036 415676 492088 415682
rect 492036 415618 492088 415624
rect 512736 415676 512788 415682
rect 512736 415618 512788 415624
rect 492048 413916 492076 415618
rect 501696 415608 501748 415614
rect 501696 415550 501748 415556
rect 501708 413916 501736 415550
rect 511448 415540 511500 415546
rect 511448 415482 511500 415488
rect 511356 415472 511408 415478
rect 511356 415414 511408 415420
rect 511368 413916 511396 415414
rect 491668 395072 491720 395078
rect 491668 395014 491720 395020
rect 491680 394754 491708 395014
rect 511460 394754 511488 415482
rect 512644 415472 512696 415478
rect 512644 415414 512696 415420
rect 491680 394726 492062 394754
rect 511382 394726 511488 394754
rect 501708 391814 501736 394060
rect 512656 391814 512684 415414
rect 512748 395078 512776 415618
rect 529664 415540 529716 415546
rect 529664 415482 529716 415488
rect 529676 413916 529704 415482
rect 539324 415472 539376 415478
rect 539324 415414 539376 415420
rect 540244 415472 540296 415478
rect 540244 415414 540296 415420
rect 539336 413916 539364 415414
rect 519004 413222 520030 413250
rect 518806 404288 518862 404297
rect 518806 404223 518862 404232
rect 513378 403608 513434 403617
rect 513378 403543 513434 403552
rect 512736 395072 512788 395078
rect 512736 395014 512788 395020
rect 513392 394602 513420 403543
rect 518820 394602 518848 404223
rect 513380 394596 513432 394602
rect 513380 394538 513432 394544
rect 518808 394596 518860 394602
rect 518808 394538 518860 394544
rect 519004 391814 519032 413222
rect 519636 395072 519688 395078
rect 519636 395014 519688 395020
rect 519648 394754 519676 395014
rect 519648 394726 520030 394754
rect 501696 391808 501748 391814
rect 501696 391750 501748 391756
rect 512644 391808 512696 391814
rect 512644 391750 512696 391756
rect 518992 391808 519044 391814
rect 518992 391750 519044 391756
rect 529676 391746 529704 394060
rect 539336 391950 539364 394060
rect 539324 391944 539376 391950
rect 539324 391886 539376 391892
rect 540256 391746 540284 415414
rect 529664 391740 529716 391746
rect 529664 391682 529716 391688
rect 540244 391740 540296 391746
rect 540244 391682 540296 391688
rect 492036 389428 492088 389434
rect 492036 389370 492088 389376
rect 512736 389428 512788 389434
rect 512736 389370 512788 389376
rect 492048 386852 492076 389370
rect 501696 389360 501748 389366
rect 501696 389302 501748 389308
rect 501708 386852 501736 389302
rect 511448 389292 511500 389298
rect 511448 389234 511500 389240
rect 511356 389224 511408 389230
rect 511356 389166 511408 389172
rect 511368 386852 511396 389166
rect 491668 368892 491720 368898
rect 491668 368834 491720 368840
rect 491680 367690 491708 368834
rect 511460 367690 511488 389234
rect 512644 389224 512696 389230
rect 512644 389166 512696 389172
rect 491680 367662 492062 367690
rect 511382 367662 511488 367690
rect 501708 365566 501736 367132
rect 512656 365566 512684 389166
rect 512748 368762 512776 389370
rect 529664 389292 529716 389298
rect 529664 389234 529716 389240
rect 529676 386852 529704 389234
rect 539324 389224 539376 389230
rect 539324 389166 539376 389172
rect 540244 389224 540296 389230
rect 540244 389166 540296 389172
rect 539336 386852 539364 389166
rect 519556 386294 520030 386322
rect 518806 377088 518862 377097
rect 518806 377023 518862 377032
rect 513378 376000 513434 376009
rect 513378 375935 513434 375944
rect 512736 368756 512788 368762
rect 512736 368698 512788 368704
rect 513392 368422 513420 375935
rect 518820 368422 518848 377023
rect 519556 373994 519584 386294
rect 519004 373966 519584 373994
rect 513380 368416 513432 368422
rect 513380 368358 513432 368364
rect 518808 368416 518860 368422
rect 518808 368358 518860 368364
rect 519004 365566 519032 373966
rect 519636 368756 519688 368762
rect 519636 368698 519688 368704
rect 519648 367690 519676 368698
rect 519648 367662 520030 367690
rect 501696 365560 501748 365566
rect 501696 365502 501748 365508
rect 512644 365560 512696 365566
rect 512644 365502 512696 365508
rect 518992 365560 519044 365566
rect 518992 365502 519044 365508
rect 529676 365498 529704 367132
rect 539336 365702 539364 367132
rect 539324 365696 539376 365702
rect 539324 365638 539376 365644
rect 540256 365498 540284 389166
rect 540886 376000 540942 376009
rect 540886 375935 540942 375944
rect 540900 368490 540928 375935
rect 540888 368484 540940 368490
rect 540888 368426 540940 368432
rect 529664 365492 529716 365498
rect 529664 365434 529716 365440
rect 540244 365492 540296 365498
rect 540244 365434 540296 365440
rect 492036 361820 492088 361826
rect 492036 361762 492088 361768
rect 512736 361820 512788 361826
rect 512736 361762 512788 361768
rect 492048 359924 492076 361762
rect 501696 361752 501748 361758
rect 501696 361694 501748 361700
rect 501708 359924 501736 361694
rect 511448 361684 511500 361690
rect 511448 361626 511500 361632
rect 511356 361616 511408 361622
rect 511356 361558 511408 361564
rect 511368 359924 511396 361558
rect 491668 341420 491720 341426
rect 491668 341362 491720 341368
rect 491680 340762 491708 341362
rect 511460 340762 511488 361626
rect 512644 361616 512696 361622
rect 512644 361558 512696 361564
rect 491680 340734 492062 340762
rect 511382 340734 511488 340762
rect 501708 337958 501736 340068
rect 512656 337958 512684 361558
rect 512748 341970 512776 361762
rect 529664 361684 529716 361690
rect 529664 361626 529716 361632
rect 529676 359924 529704 361626
rect 539324 361616 539376 361622
rect 539324 361558 539376 361564
rect 540244 361616 540296 361622
rect 540244 361558 540296 361564
rect 539336 359924 539364 361558
rect 519004 359230 520030 359258
rect 518806 350296 518862 350305
rect 518806 350231 518862 350240
rect 513378 349616 513434 349625
rect 513378 349551 513434 349560
rect 512736 341964 512788 341970
rect 512736 341906 512788 341912
rect 513392 340746 513420 349551
rect 518820 340814 518848 350231
rect 518808 340808 518860 340814
rect 518808 340750 518860 340756
rect 513380 340740 513432 340746
rect 513380 340682 513432 340688
rect 519004 337958 519032 359230
rect 519636 341964 519688 341970
rect 519636 341906 519688 341912
rect 519648 340762 519676 341906
rect 519648 340734 520030 340762
rect 539350 340746 539548 340762
rect 539350 340740 539560 340746
rect 539350 340734 539508 340740
rect 539508 340682 539560 340688
rect 501696 337952 501748 337958
rect 501696 337894 501748 337900
rect 512644 337952 512696 337958
rect 512644 337894 512696 337900
rect 518992 337952 519044 337958
rect 518992 337894 519044 337900
rect 529676 337890 529704 340068
rect 540256 337890 540284 361558
rect 529664 337884 529716 337890
rect 529664 337826 529716 337832
rect 540244 337884 540296 337890
rect 540244 337826 540296 337832
rect 492036 335572 492088 335578
rect 492036 335514 492088 335520
rect 512736 335572 512788 335578
rect 512736 335514 512788 335520
rect 492048 332860 492076 335514
rect 501696 335504 501748 335510
rect 501696 335446 501748 335452
rect 501708 332860 501736 335446
rect 511448 335436 511500 335442
rect 511448 335378 511500 335384
rect 511356 335368 511408 335374
rect 511356 335310 511408 335316
rect 511368 332860 511396 335310
rect 491668 315988 491720 315994
rect 491668 315930 491720 315936
rect 491680 313698 491708 315930
rect 511460 313698 511488 335378
rect 512644 335368 512696 335374
rect 512644 335310 512696 335316
rect 491680 313670 492062 313698
rect 511382 313670 511488 313698
rect 501708 311710 501736 313140
rect 512656 311710 512684 335310
rect 512748 315314 512776 335514
rect 529664 335436 529716 335442
rect 529664 335378 529716 335384
rect 529676 332860 529704 335378
rect 539324 335368 539376 335374
rect 539324 335310 539376 335316
rect 540244 335368 540296 335374
rect 540244 335310 540296 335316
rect 539336 332860 539364 335310
rect 519004 332302 520030 332330
rect 513380 331288 513432 331294
rect 513380 331230 513432 331236
rect 513392 322833 513420 331230
rect 518806 322960 518862 322969
rect 518806 322895 518862 322904
rect 513378 322824 513434 322833
rect 513378 322759 513434 322768
rect 512736 315308 512788 315314
rect 512736 315250 512788 315256
rect 518820 314566 518848 322895
rect 518808 314560 518860 314566
rect 518808 314502 518860 314508
rect 519004 311710 519032 332302
rect 519636 315308 519688 315314
rect 519636 315250 519688 315256
rect 519648 313698 519676 315250
rect 519648 313670 520030 313698
rect 501696 311704 501748 311710
rect 501696 311646 501748 311652
rect 512644 311704 512696 311710
rect 512644 311646 512696 311652
rect 518992 311704 519044 311710
rect 518992 311646 519044 311652
rect 529676 311642 529704 313140
rect 539336 311846 539364 313140
rect 539324 311840 539376 311846
rect 539324 311782 539376 311788
rect 540256 311642 540284 335310
rect 529664 311636 529716 311642
rect 529664 311578 529716 311584
rect 540244 311636 540296 311642
rect 540244 311578 540296 311584
rect 492036 308032 492088 308038
rect 492036 307974 492088 307980
rect 512736 308032 512788 308038
rect 512736 307974 512788 307980
rect 492048 305932 492076 307974
rect 501696 307964 501748 307970
rect 501696 307906 501748 307912
rect 501708 305932 501736 307906
rect 511448 307896 511500 307902
rect 511448 307838 511500 307844
rect 511356 307828 511408 307834
rect 511356 307770 511408 307776
rect 511368 305932 511396 307770
rect 491668 287428 491720 287434
rect 491668 287370 491720 287376
rect 491680 286770 491708 287370
rect 511460 286770 511488 307838
rect 512644 307828 512696 307834
rect 512644 307770 512696 307776
rect 491680 286742 492062 286770
rect 511382 286742 511488 286770
rect 501708 284170 501736 286076
rect 512656 284170 512684 307770
rect 512748 287570 512776 307974
rect 529664 307896 529716 307902
rect 529664 307838 529716 307844
rect 529676 305932 529704 307838
rect 539324 307828 539376 307834
rect 539324 307770 539376 307776
rect 540244 307828 540296 307834
rect 540244 307770 540296 307776
rect 539336 305932 539364 307770
rect 519004 305238 520030 305266
rect 518806 296304 518862 296313
rect 518806 296239 518862 296248
rect 513378 295624 513434 295633
rect 513378 295559 513434 295568
rect 512736 287564 512788 287570
rect 512736 287506 512788 287512
rect 513392 286890 513420 295559
rect 518820 286958 518848 296239
rect 518808 286952 518860 286958
rect 518808 286894 518860 286900
rect 513380 286884 513432 286890
rect 513380 286826 513432 286832
rect 519004 284170 519032 305238
rect 519636 287564 519688 287570
rect 519636 287506 519688 287512
rect 519648 286770 519676 287506
rect 539508 286816 539560 286822
rect 519648 286742 520030 286770
rect 539350 286764 539508 286770
rect 539350 286758 539560 286764
rect 539350 286742 539548 286758
rect 501696 284164 501748 284170
rect 501696 284106 501748 284112
rect 512644 284164 512696 284170
rect 512644 284106 512696 284112
rect 518992 284164 519044 284170
rect 518992 284106 519044 284112
rect 529676 284102 529704 286076
rect 540256 284102 540284 307770
rect 529664 284096 529716 284102
rect 529664 284038 529716 284044
rect 540244 284096 540296 284102
rect 540244 284038 540296 284044
rect 492036 280424 492088 280430
rect 492036 280366 492088 280372
rect 512736 280424 512788 280430
rect 512736 280366 512788 280372
rect 492048 278868 492076 280366
rect 501696 280356 501748 280362
rect 501696 280298 501748 280304
rect 501708 278868 501736 280298
rect 511448 280288 511500 280294
rect 511448 280230 511500 280236
rect 511356 280220 511408 280226
rect 511356 280162 511408 280168
rect 511368 278868 511396 280162
rect 491668 262200 491720 262206
rect 491668 262142 491720 262148
rect 491680 259706 491708 262142
rect 511460 259706 511488 280230
rect 512644 280220 512696 280226
rect 512644 280162 512696 280168
rect 491680 259678 492062 259706
rect 511382 259678 511488 259706
rect 501708 256562 501736 259148
rect 512656 256562 512684 280162
rect 512748 262206 512776 280366
rect 529664 280288 529716 280294
rect 529664 280230 529716 280236
rect 529676 278868 529704 280230
rect 539324 280220 539376 280226
rect 539324 280162 539376 280168
rect 540244 280220 540296 280226
rect 540244 280162 540296 280168
rect 539336 278868 539364 280162
rect 519004 278310 520030 278338
rect 513380 277568 513432 277574
rect 513380 277510 513432 277516
rect 513392 268569 513420 277510
rect 518808 277500 518860 277506
rect 518808 277442 518860 277448
rect 518820 269249 518848 277442
rect 518806 269240 518862 269249
rect 518806 269175 518862 269184
rect 513378 268560 513434 268569
rect 513378 268495 513434 268504
rect 512736 262200 512788 262206
rect 512736 262142 512788 262148
rect 519004 256562 519032 278310
rect 519636 262200 519688 262206
rect 519636 262142 519688 262148
rect 519648 259706 519676 262142
rect 519648 259678 520030 259706
rect 501696 256556 501748 256562
rect 501696 256498 501748 256504
rect 512644 256556 512696 256562
rect 512644 256498 512696 256504
rect 518992 256556 519044 256562
rect 518992 256498 519044 256504
rect 529676 256494 529704 259148
rect 539336 256698 539364 259148
rect 539324 256692 539376 256698
rect 539324 256634 539376 256640
rect 540256 256494 540284 280162
rect 529664 256488 529716 256494
rect 529664 256430 529716 256436
rect 540244 256488 540296 256494
rect 540244 256430 540296 256436
rect 492036 254176 492088 254182
rect 492036 254118 492088 254124
rect 512736 254176 512788 254182
rect 512736 254118 512788 254124
rect 492048 251940 492076 254118
rect 501696 254108 501748 254114
rect 501696 254050 501748 254056
rect 501708 251940 501736 254050
rect 511448 254040 511500 254046
rect 511448 253982 511500 253988
rect 511356 253972 511408 253978
rect 511356 253914 511408 253920
rect 511368 251940 511396 253914
rect 491668 233436 491720 233442
rect 491668 233378 491720 233384
rect 491680 232778 491708 233378
rect 511460 232778 511488 253982
rect 512644 253972 512696 253978
rect 512644 253914 512696 253920
rect 491680 232750 492062 232778
rect 511382 232750 511488 232778
rect 501708 230314 501736 232084
rect 512656 230314 512684 253914
rect 512748 234258 512776 254118
rect 529664 254040 529716 254046
rect 529664 253982 529716 253988
rect 529676 251940 529704 253982
rect 539324 253972 539376 253978
rect 539324 253914 539376 253920
rect 540244 253972 540296 253978
rect 540244 253914 540296 253920
rect 539336 251940 539364 253914
rect 519004 251246 520030 251274
rect 518806 242312 518862 242321
rect 518806 242247 518862 242256
rect 513378 241632 513434 241641
rect 513378 241567 513434 241576
rect 512736 234252 512788 234258
rect 512736 234194 512788 234200
rect 513392 233238 513420 241567
rect 518820 233238 518848 242247
rect 513380 233232 513432 233238
rect 513380 233174 513432 233180
rect 518808 233232 518860 233238
rect 518808 233174 518860 233180
rect 519004 230314 519032 251246
rect 519636 234252 519688 234258
rect 519636 234194 519688 234200
rect 519648 232778 519676 234194
rect 539508 233164 539560 233170
rect 539508 233106 539560 233112
rect 539520 232778 539548 233106
rect 519648 232750 520030 232778
rect 539350 232750 539548 232778
rect 501696 230308 501748 230314
rect 501696 230250 501748 230256
rect 512644 230308 512696 230314
rect 512644 230250 512696 230256
rect 518992 230308 519044 230314
rect 518992 230250 519044 230256
rect 529676 230246 529704 232084
rect 540256 230246 540284 253914
rect 529664 230240 529716 230246
rect 529664 230182 529716 230188
rect 540244 230240 540296 230246
rect 540244 230182 540296 230188
rect 492036 226568 492088 226574
rect 492036 226510 492088 226516
rect 512736 226568 512788 226574
rect 512736 226510 512788 226516
rect 492048 224876 492076 226510
rect 501696 226500 501748 226506
rect 501696 226442 501748 226448
rect 501708 224876 501736 226442
rect 511448 226432 511500 226438
rect 511448 226374 511500 226380
rect 511356 226364 511408 226370
rect 511356 226306 511408 226312
rect 511368 224876 511396 226306
rect 491668 207460 491720 207466
rect 491668 207402 491720 207408
rect 491680 205714 491708 207402
rect 511460 205714 511488 226374
rect 512644 226364 512696 226370
rect 512644 226306 512696 226312
rect 491680 205686 492062 205714
rect 511382 205686 511488 205714
rect 501708 202706 501736 205020
rect 512656 202706 512684 226306
rect 512748 207330 512776 226510
rect 529664 226432 529716 226438
rect 529664 226374 529716 226380
rect 529676 224876 529704 226374
rect 539324 226364 539376 226370
rect 539324 226306 539376 226312
rect 540244 226364 540296 226370
rect 540244 226306 540296 226312
rect 539336 224876 539364 226306
rect 519004 224318 520030 224346
rect 518806 215248 518862 215257
rect 518806 215183 518862 215192
rect 513378 214568 513434 214577
rect 513378 214503 513434 214512
rect 512736 207324 512788 207330
rect 512736 207266 512788 207272
rect 513392 205494 513420 214503
rect 518820 205562 518848 215183
rect 518808 205556 518860 205562
rect 518808 205498 518860 205504
rect 513380 205488 513432 205494
rect 513380 205430 513432 205436
rect 519004 202706 519032 224318
rect 519636 207324 519688 207330
rect 519636 207266 519688 207272
rect 519648 205714 519676 207266
rect 519648 205686 520030 205714
rect 539508 205488 539560 205494
rect 539350 205436 539508 205442
rect 539350 205430 539560 205436
rect 539350 205414 539548 205430
rect 501696 202700 501748 202706
rect 501696 202642 501748 202648
rect 512644 202700 512696 202706
rect 512644 202642 512696 202648
rect 518992 202700 519044 202706
rect 518992 202642 519044 202648
rect 529676 202638 529704 205020
rect 540256 202638 540284 226306
rect 529664 202632 529716 202638
rect 529664 202574 529716 202580
rect 540244 202632 540296 202638
rect 540244 202574 540296 202580
rect 492036 200388 492088 200394
rect 492036 200330 492088 200336
rect 512736 200388 512788 200394
rect 512736 200330 512788 200336
rect 492048 197948 492076 200330
rect 501696 200320 501748 200326
rect 501696 200262 501748 200268
rect 501708 197948 501736 200262
rect 511448 200252 511500 200258
rect 511448 200194 511500 200200
rect 511356 200184 511408 200190
rect 511356 200126 511408 200132
rect 511368 197948 511396 200126
rect 491668 179716 491720 179722
rect 491668 179658 491720 179664
rect 491680 178786 491708 179658
rect 511460 178786 511488 200194
rect 512644 200184 512696 200190
rect 512644 200126 512696 200132
rect 491680 178758 492062 178786
rect 511382 178758 511488 178786
rect 501708 176526 501736 178092
rect 512656 176526 512684 200126
rect 512748 179858 512776 200330
rect 529664 200252 529716 200258
rect 529664 200194 529716 200200
rect 529676 197948 529704 200194
rect 539324 200184 539376 200190
rect 539324 200126 539376 200132
rect 540244 200184 540296 200190
rect 540244 200126 540296 200132
rect 539336 197948 539364 200126
rect 519004 197254 520030 197282
rect 518806 188320 518862 188329
rect 518806 188255 518862 188264
rect 513378 187640 513434 187649
rect 513378 187575 513434 187584
rect 512736 179852 512788 179858
rect 512736 179794 512788 179800
rect 513392 179246 513420 187575
rect 518820 179314 518848 188255
rect 518808 179308 518860 179314
rect 518808 179250 518860 179256
rect 513380 179240 513432 179246
rect 513380 179182 513432 179188
rect 519004 176526 519032 197254
rect 519636 179852 519688 179858
rect 519636 179794 519688 179800
rect 519648 178786 519676 179794
rect 519648 178758 520030 178786
rect 501696 176520 501748 176526
rect 501696 176462 501748 176468
rect 512644 176520 512696 176526
rect 512644 176462 512696 176468
rect 518992 176520 519044 176526
rect 518992 176462 519044 176468
rect 529676 176458 529704 178092
rect 539336 176662 539364 178092
rect 539324 176656 539376 176662
rect 539324 176598 539376 176604
rect 540256 176458 540284 200126
rect 529664 176452 529716 176458
rect 529664 176394 529716 176400
rect 540244 176452 540296 176458
rect 540244 176394 540296 176400
rect 492036 172780 492088 172786
rect 492036 172722 492088 172728
rect 512736 172780 512788 172786
rect 512736 172722 512788 172728
rect 492048 170884 492076 172722
rect 501696 172712 501748 172718
rect 501696 172654 501748 172660
rect 501708 170884 501736 172654
rect 511448 172644 511500 172650
rect 511448 172586 511500 172592
rect 511356 172576 511408 172582
rect 511356 172518 511408 172524
rect 511368 170884 511396 172518
rect 491668 152516 491720 152522
rect 491668 152458 491720 152464
rect 491680 151722 491708 152458
rect 511460 151722 511488 172586
rect 512644 172576 512696 172582
rect 512644 172518 512696 172524
rect 491680 151694 492062 151722
rect 511382 151694 511488 151722
rect 501708 148918 501736 151028
rect 512656 148918 512684 172518
rect 512748 152250 512776 172722
rect 529664 172644 529716 172650
rect 529664 172586 529716 172592
rect 529676 170884 529704 172586
rect 539324 172576 539376 172582
rect 539324 172518 539376 172524
rect 540244 172576 540296 172582
rect 540244 172518 540296 172524
rect 539336 170884 539364 172518
rect 519004 170326 520030 170354
rect 518806 161256 518862 161265
rect 518806 161191 518862 161200
rect 513378 160576 513434 160585
rect 513378 160511 513434 160520
rect 512736 152244 512788 152250
rect 512736 152186 512788 152192
rect 513392 151638 513420 160511
rect 518820 151706 518848 161191
rect 518808 151700 518860 151706
rect 518808 151642 518860 151648
rect 513380 151632 513432 151638
rect 513380 151574 513432 151580
rect 519004 148918 519032 170326
rect 519636 152244 519688 152250
rect 519636 152186 519688 152192
rect 519648 151722 519676 152186
rect 519648 151694 520030 151722
rect 539508 151632 539560 151638
rect 539350 151580 539508 151586
rect 539350 151574 539560 151580
rect 539350 151558 539548 151574
rect 501696 148912 501748 148918
rect 501696 148854 501748 148860
rect 512644 148912 512696 148918
rect 512644 148854 512696 148860
rect 518992 148912 519044 148918
rect 518992 148854 519044 148860
rect 529676 148850 529704 151028
rect 540256 148850 540284 172518
rect 529664 148844 529716 148850
rect 529664 148786 529716 148792
rect 540244 148844 540296 148850
rect 540244 148786 540296 148792
rect 492036 146532 492088 146538
rect 492036 146474 492088 146480
rect 512736 146532 512788 146538
rect 512736 146474 512788 146480
rect 492048 143956 492076 146474
rect 501696 146464 501748 146470
rect 501696 146406 501748 146412
rect 501708 143956 501736 146406
rect 511448 146396 511500 146402
rect 511448 146338 511500 146344
rect 511356 146328 511408 146334
rect 511356 146270 511408 146276
rect 511368 143956 511396 146270
rect 491668 126948 491720 126954
rect 491668 126890 491720 126896
rect 491680 124794 491708 126890
rect 511460 124794 511488 146338
rect 512644 146328 512696 146334
rect 512644 146270 512696 146276
rect 491680 124766 492062 124794
rect 511382 124766 511488 124794
rect 501708 122670 501736 124100
rect 512656 122670 512684 146270
rect 512748 126954 512776 146474
rect 529664 146396 529716 146402
rect 529664 146338 529716 146344
rect 529676 143956 529704 146338
rect 539324 146328 539376 146334
rect 539324 146270 539376 146276
rect 540244 146328 540296 146334
rect 540244 146270 540296 146276
rect 539336 143956 539364 146270
rect 519004 143262 520030 143290
rect 518806 134328 518862 134337
rect 518806 134263 518862 134272
rect 513378 133648 513434 133657
rect 513378 133583 513434 133592
rect 512736 126948 512788 126954
rect 512736 126890 512788 126896
rect 513392 125458 513420 133583
rect 518820 125526 518848 134263
rect 518808 125520 518860 125526
rect 518808 125462 518860 125468
rect 513380 125452 513432 125458
rect 513380 125394 513432 125400
rect 519004 122670 519032 143262
rect 519636 126948 519688 126954
rect 519636 126890 519688 126896
rect 519648 124794 519676 126890
rect 519648 124766 520030 124794
rect 501696 122664 501748 122670
rect 501696 122606 501748 122612
rect 512644 122664 512696 122670
rect 512644 122606 512696 122612
rect 518992 122664 519044 122670
rect 518992 122606 519044 122612
rect 529676 122602 529704 124100
rect 539336 122806 539364 124100
rect 539324 122800 539376 122806
rect 539324 122742 539376 122748
rect 540256 122602 540284 146270
rect 529664 122596 529716 122602
rect 529664 122538 529716 122544
rect 540244 122596 540296 122602
rect 540244 122538 540296 122544
rect 492036 118924 492088 118930
rect 492036 118866 492088 118872
rect 512736 118924 512788 118930
rect 512736 118866 512788 118872
rect 492048 116892 492076 118866
rect 501696 118856 501748 118862
rect 501696 118798 501748 118804
rect 501708 116892 501736 118798
rect 511448 118788 511500 118794
rect 511448 118730 511500 118736
rect 511356 118720 511408 118726
rect 511356 118662 511408 118668
rect 511368 116892 511396 118662
rect 491668 98660 491720 98666
rect 491668 98602 491720 98608
rect 491680 97730 491708 98602
rect 511460 97730 511488 118730
rect 512644 118720 512696 118726
rect 512644 118662 512696 118668
rect 491680 97702 492062 97730
rect 511382 97702 511488 97730
rect 501708 95062 501736 97036
rect 512656 95062 512684 118662
rect 512748 98598 512776 118866
rect 529664 118788 529716 118794
rect 529664 118730 529716 118736
rect 529676 116892 529704 118730
rect 539324 118720 539376 118726
rect 539324 118662 539376 118668
rect 540244 118720 540296 118726
rect 540244 118662 540296 118668
rect 539336 116892 539364 118662
rect 519004 116334 520030 116362
rect 518806 107264 518862 107273
rect 518806 107199 518862 107208
rect 513378 106584 513434 106593
rect 513378 106519 513434 106528
rect 512736 98592 512788 98598
rect 512736 98534 512788 98540
rect 513392 97918 513420 106519
rect 518820 97918 518848 107199
rect 513380 97912 513432 97918
rect 513380 97854 513432 97860
rect 518808 97912 518860 97918
rect 518808 97854 518860 97860
rect 519004 95062 519032 116334
rect 519636 98592 519688 98598
rect 519636 98534 519688 98540
rect 519648 97730 519676 98534
rect 539508 97844 539560 97850
rect 539508 97786 539560 97792
rect 539520 97730 539548 97786
rect 519648 97702 520030 97730
rect 539350 97702 539548 97730
rect 501696 95056 501748 95062
rect 501696 94998 501748 95004
rect 512644 95056 512696 95062
rect 512644 94998 512696 95004
rect 518992 95056 519044 95062
rect 518992 94998 519044 95004
rect 529676 94994 529704 97036
rect 540256 94994 540284 118662
rect 529664 94988 529716 94994
rect 529664 94930 529716 94936
rect 540244 94988 540296 94994
rect 540244 94930 540296 94936
rect 501696 91248 501748 91254
rect 501696 91190 501748 91196
rect 511448 91248 511500 91254
rect 511448 91190 511500 91196
rect 529664 91248 529716 91254
rect 529664 91190 529716 91196
rect 492036 91180 492088 91186
rect 492036 91122 492088 91128
rect 492048 89964 492076 91122
rect 501708 89964 501736 91190
rect 511356 91112 511408 91118
rect 511356 91054 511408 91060
rect 511368 89964 511396 91054
rect 491668 72276 491720 72282
rect 491668 72218 491720 72224
rect 491680 70666 491708 72218
rect 511460 70666 511488 91190
rect 512736 91180 512788 91186
rect 512736 91122 512788 91128
rect 512644 91112 512696 91118
rect 512644 91054 512696 91060
rect 491680 70638 492062 70666
rect 511382 70638 511488 70666
rect 501708 68882 501736 70108
rect 512656 68882 512684 91054
rect 512748 72146 512776 91122
rect 529676 89964 529704 91190
rect 539324 91112 539376 91118
rect 539324 91054 539376 91060
rect 540244 91112 540296 91118
rect 540244 91054 540296 91060
rect 539336 89964 539364 91054
rect 519004 89270 520030 89298
rect 518808 88392 518860 88398
rect 518808 88334 518860 88340
rect 518820 80345 518848 88334
rect 518806 80336 518862 80345
rect 518806 80271 518862 80280
rect 513378 79656 513434 79665
rect 513378 79591 513434 79600
rect 512736 72140 512788 72146
rect 512736 72082 512788 72088
rect 513392 71670 513420 79591
rect 513380 71664 513432 71670
rect 513380 71606 513432 71612
rect 519004 68882 519032 89270
rect 519636 72140 519688 72146
rect 519636 72082 519688 72088
rect 519648 70666 519676 72082
rect 519648 70638 520030 70666
rect 501696 68876 501748 68882
rect 501696 68818 501748 68824
rect 512644 68876 512696 68882
rect 512644 68818 512696 68824
rect 518992 68876 519044 68882
rect 518992 68818 519044 68824
rect 529676 68814 529704 70108
rect 539336 69018 539364 70108
rect 539324 69012 539376 69018
rect 539324 68954 539376 68960
rect 540256 68814 540284 91054
rect 529664 68808 529716 68814
rect 529664 68750 529716 68756
rect 540244 68808 540296 68814
rect 540244 68750 540296 68756
rect 501696 65068 501748 65074
rect 501696 65010 501748 65016
rect 511448 65068 511500 65074
rect 511448 65010 511500 65016
rect 529664 65068 529716 65074
rect 529664 65010 529716 65016
rect 492036 65000 492088 65006
rect 492036 64942 492088 64948
rect 492048 62900 492076 64942
rect 501708 62900 501736 65010
rect 511356 64932 511408 64938
rect 511356 64874 511408 64880
rect 511368 62900 511396 64874
rect 491668 44668 491720 44674
rect 491668 44610 491720 44616
rect 491680 43738 491708 44610
rect 511460 43738 511488 65010
rect 512736 65000 512788 65006
rect 512736 64942 512788 64948
rect 512644 64932 512696 64938
rect 512644 64874 512696 64880
rect 491680 43710 492062 43738
rect 511382 43710 511488 43738
rect 501708 41274 501736 43044
rect 512656 41274 512684 64874
rect 512748 44742 512776 64942
rect 529676 62900 529704 65010
rect 539324 64932 539376 64938
rect 539324 64874 539376 64880
rect 540244 64932 540296 64938
rect 540244 64874 540296 64880
rect 539336 62900 539364 64874
rect 519004 62206 520030 62234
rect 518806 53272 518862 53281
rect 518806 53207 518862 53216
rect 513378 52592 513434 52601
rect 513378 52527 513434 52536
rect 512736 44736 512788 44742
rect 512736 44678 512788 44684
rect 513392 44130 513420 52527
rect 518820 44130 518848 53207
rect 513380 44124 513432 44130
rect 513380 44066 513432 44072
rect 518808 44124 518860 44130
rect 518808 44066 518860 44072
rect 519004 41274 519032 62206
rect 519636 44736 519688 44742
rect 519636 44678 519688 44684
rect 519648 43738 519676 44678
rect 539508 44056 539560 44062
rect 539508 43998 539560 44004
rect 539520 43738 539548 43998
rect 519648 43710 520030 43738
rect 539350 43710 539548 43738
rect 501696 41268 501748 41274
rect 501696 41210 501748 41216
rect 512644 41268 512696 41274
rect 512644 41210 512696 41216
rect 518992 41268 519044 41274
rect 518992 41210 519044 41216
rect 529676 41206 529704 43044
rect 540256 41206 540284 64874
rect 529664 41200 529716 41206
rect 529664 41142 529716 41148
rect 540244 41200 540296 41206
rect 540244 41142 540296 41148
rect 501696 37460 501748 37466
rect 501696 37402 501748 37408
rect 492036 37392 492088 37398
rect 492036 37334 492088 37340
rect 492048 35972 492076 37334
rect 501708 35972 501736 37402
rect 512736 37392 512788 37398
rect 512736 37334 512788 37340
rect 518164 37392 518216 37398
rect 518164 37334 518216 37340
rect 529664 37392 529716 37398
rect 529664 37334 529716 37340
rect 511356 37324 511408 37330
rect 511356 37266 511408 37272
rect 512644 37324 512696 37330
rect 512644 37266 512696 37272
rect 511368 35972 511396 37266
rect 491668 18012 491720 18018
rect 491668 17954 491720 17960
rect 491680 16674 491708 17954
rect 491680 16646 492062 16674
rect 501708 13598 501736 16116
rect 511368 13802 511396 16116
rect 511356 13796 511408 13802
rect 511356 13738 511408 13744
rect 512656 13598 512684 37266
rect 512748 18018 512776 37334
rect 513380 34604 513432 34610
rect 513380 34546 513432 34552
rect 513392 25673 513420 34546
rect 513378 25664 513434 25673
rect 513378 25599 513434 25608
rect 512736 18012 512788 18018
rect 512736 17954 512788 17960
rect 518176 13802 518204 37334
rect 529676 35972 529704 37334
rect 539324 37324 539376 37330
rect 539324 37266 539376 37272
rect 539336 35972 539364 37266
rect 519004 35278 520030 35306
rect 518808 34604 518860 34610
rect 518808 34546 518860 34552
rect 518820 26353 518848 34546
rect 518806 26344 518862 26353
rect 518806 26279 518862 26288
rect 518164 13796 518216 13802
rect 518164 13738 518216 13744
rect 519004 13598 519032 35278
rect 519636 18012 519688 18018
rect 519636 17954 519688 17960
rect 519648 16674 519676 17954
rect 519648 16646 520030 16674
rect 539508 16584 539560 16590
rect 539350 16532 539508 16538
rect 539350 16526 539560 16532
rect 539350 16510 539548 16526
rect 490564 13592 490616 13598
rect 490564 13534 490616 13540
rect 501696 13592 501748 13598
rect 501696 13534 501748 13540
rect 512644 13592 512696 13598
rect 512644 13534 512696 13540
rect 518992 13592 519044 13598
rect 518992 13534 519044 13540
rect 529676 13462 529704 16116
rect 64144 13456 64196 13462
rect 64144 13398 64196 13404
rect 72056 13456 72108 13462
rect 72056 13398 72108 13404
rect 99472 13456 99524 13462
rect 99472 13398 99524 13404
rect 127072 13456 127124 13462
rect 127072 13398 127124 13404
rect 238852 13456 238904 13462
rect 238852 13398 238904 13404
rect 268016 13456 268068 13462
rect 268016 13398 268068 13404
rect 323032 13456 323084 13462
rect 323032 13398 323084 13404
rect 352012 13456 352064 13462
rect 352012 13398 352064 13404
rect 379612 13456 379664 13462
rect 379612 13398 379664 13404
rect 408040 13456 408092 13462
rect 408040 13398 408092 13404
rect 434812 13456 434864 13462
rect 434812 13398 434864 13404
rect 463700 13456 463752 13462
rect 463700 13398 463752 13404
rect 529664 13456 529716 13462
rect 529664 13398 529716 13404
rect 541636 13326 541664 673814
rect 542372 673577 542400 683130
rect 542358 673568 542414 673577
rect 542358 673503 542414 673512
rect 543016 662318 543044 685918
rect 557552 683754 557580 685918
rect 567200 685908 567252 685914
rect 567200 685850 567252 685856
rect 567212 683754 567240 685850
rect 557552 683726 557704 683754
rect 567212 683726 567364 683754
rect 545118 674248 545174 674257
rect 545118 674183 545174 674192
rect 545132 673878 545160 674183
rect 545120 673872 545172 673878
rect 545120 673814 545172 673820
rect 569958 673568 570014 673577
rect 569958 673503 570014 673512
rect 567844 670744 567896 670750
rect 567844 670686 567896 670692
rect 547892 664006 548044 664034
rect 547892 662386 547920 664006
rect 547880 662380 547932 662386
rect 547880 662322 547932 662328
rect 543004 662312 543056 662318
rect 543004 662254 543056 662260
rect 547880 658980 547932 658986
rect 547880 658922 547932 658928
rect 543004 658368 543056 658374
rect 543004 658310 543056 658316
rect 542360 655580 542412 655586
rect 542360 655522 542412 655528
rect 542372 646649 542400 655522
rect 542358 646640 542414 646649
rect 542358 646575 542414 646584
rect 543016 634778 543044 658310
rect 545764 657552 545816 657558
rect 545764 657494 545816 657500
rect 545776 647329 545804 657494
rect 547892 656826 547920 658922
rect 557540 658368 557592 658374
rect 557540 658310 557592 658316
rect 557552 656826 557580 658310
rect 567200 658300 567252 658306
rect 567200 658242 567252 658248
rect 567212 656826 567240 658242
rect 547892 656798 548044 656826
rect 557552 656798 557704 656826
rect 567212 656798 567364 656826
rect 545762 647320 545818 647329
rect 545762 647255 545818 647264
rect 547892 637078 548044 637106
rect 557552 637078 557704 637106
rect 567212 637078 567364 637106
rect 543004 634772 543056 634778
rect 543004 634714 543056 634720
rect 547892 634642 547920 637078
rect 547880 634636 547932 634642
rect 547880 634578 547932 634584
rect 557552 634506 557580 637078
rect 567212 634710 567240 637078
rect 567200 634704 567252 634710
rect 567200 634646 567252 634652
rect 557540 634500 557592 634506
rect 557540 634442 557592 634448
rect 547880 632732 547932 632738
rect 547880 632674 547932 632680
rect 543004 632188 543056 632194
rect 543004 632130 543056 632136
rect 542358 619576 542414 619585
rect 542358 619511 542414 619520
rect 542372 611318 542400 619511
rect 542360 611312 542412 611318
rect 542360 611254 542412 611260
rect 543016 608598 543044 632130
rect 545764 629944 545816 629950
rect 545764 629886 545816 629892
rect 545776 620265 545804 629886
rect 547892 629762 547920 632674
rect 557540 632188 557592 632194
rect 557540 632130 557592 632136
rect 557552 629762 557580 632130
rect 567200 632120 567252 632126
rect 567200 632062 567252 632068
rect 567212 629762 567240 632062
rect 547892 629734 548044 629762
rect 557552 629734 557704 629762
rect 567212 629734 567364 629762
rect 545762 620256 545818 620265
rect 545762 620191 545818 620200
rect 547892 610014 548044 610042
rect 557552 610014 557704 610042
rect 567212 610014 567364 610042
rect 543004 608592 543056 608598
rect 543004 608534 543056 608540
rect 547892 608462 547920 610014
rect 547880 608456 547932 608462
rect 547880 608398 547932 608404
rect 557552 608326 557580 610014
rect 567212 608530 567240 610014
rect 567200 608524 567252 608530
rect 567200 608466 567252 608472
rect 557540 608320 557592 608326
rect 557540 608262 557592 608268
rect 547880 605124 547932 605130
rect 547880 605066 547932 605072
rect 543004 604580 543056 604586
rect 543004 604522 543056 604528
rect 542358 592648 542414 592657
rect 542358 592583 542414 592592
rect 542372 583710 542400 592583
rect 542360 583704 542412 583710
rect 542360 583646 542412 583652
rect 543016 583574 543044 604522
rect 547892 602834 547920 605066
rect 557540 604580 557592 604586
rect 557540 604522 557592 604528
rect 557552 602834 557580 604522
rect 567200 604512 567252 604518
rect 567200 604454 567252 604460
rect 567212 602834 567240 604454
rect 547892 602806 548044 602834
rect 557552 602806 557704 602834
rect 567212 602806 567364 602834
rect 545764 602404 545816 602410
rect 545764 602346 545816 602352
rect 545776 593337 545804 602346
rect 545762 593328 545818 593337
rect 545762 593263 545818 593272
rect 543004 583568 543056 583574
rect 543004 583510 543056 583516
rect 547892 583086 548044 583114
rect 557552 583086 557704 583114
rect 567212 583086 567364 583114
rect 547892 580854 547920 583086
rect 547880 580848 547932 580854
rect 547880 580790 547932 580796
rect 557552 580718 557580 583086
rect 567212 580922 567240 583086
rect 567200 580916 567252 580922
rect 567200 580858 567252 580864
rect 557540 580712 557592 580718
rect 557540 580654 557592 580660
rect 547880 578944 547932 578950
rect 547880 578886 547932 578892
rect 543004 578332 543056 578338
rect 543004 578274 543056 578280
rect 542358 565584 542414 565593
rect 542358 565519 542414 565528
rect 542372 557530 542400 565519
rect 542360 557524 542412 557530
rect 542360 557466 542412 557472
rect 543016 554742 543044 578274
rect 545764 576156 545816 576162
rect 545764 576098 545816 576104
rect 545776 566273 545804 576098
rect 547892 575906 547920 578886
rect 557540 578332 557592 578338
rect 557540 578274 557592 578280
rect 557552 575906 557580 578274
rect 567200 578264 567252 578270
rect 567200 578206 567252 578212
rect 567212 575906 567240 578206
rect 547892 575878 548044 575906
rect 557552 575878 557704 575906
rect 567212 575878 567364 575906
rect 545762 566264 545818 566273
rect 545762 566199 545818 566208
rect 547892 556022 548044 556050
rect 557552 556022 557704 556050
rect 567212 556022 567364 556050
rect 543004 554736 543056 554742
rect 543004 554678 543056 554684
rect 547892 554606 547920 556022
rect 547880 554600 547932 554606
rect 547880 554542 547932 554548
rect 557552 554470 557580 556022
rect 567212 554674 567240 556022
rect 567200 554668 567252 554674
rect 567200 554610 567252 554616
rect 557540 554464 557592 554470
rect 557540 554406 557592 554412
rect 547880 551336 547932 551342
rect 547880 551278 547932 551284
rect 543004 550724 543056 550730
rect 543004 550666 543056 550672
rect 542358 538656 542414 538665
rect 542358 538591 542414 538600
rect 542372 529922 542400 538591
rect 542360 529916 542412 529922
rect 542360 529858 542412 529864
rect 543016 527134 543044 550666
rect 547892 548842 547920 551278
rect 557540 550724 557592 550730
rect 557540 550666 557592 550672
rect 557552 548842 557580 550666
rect 567200 550656 567252 550662
rect 567200 550598 567252 550604
rect 567212 548842 567240 550598
rect 547892 548814 548044 548842
rect 557552 548814 557704 548842
rect 567212 548814 567364 548842
rect 545764 548548 545816 548554
rect 545764 548490 545816 548496
rect 545776 539345 545804 548490
rect 545762 539336 545818 539345
rect 545762 539271 545818 539280
rect 547892 529094 548044 529122
rect 557552 529094 557704 529122
rect 567212 529094 567364 529122
rect 543004 527128 543056 527134
rect 543004 527070 543056 527076
rect 547892 526998 547920 529094
rect 547880 526992 547932 526998
rect 547880 526934 547932 526940
rect 557552 526862 557580 529094
rect 567212 527066 567240 529094
rect 567200 527060 567252 527066
rect 567200 527002 567252 527008
rect 557540 526856 557592 526862
rect 557540 526798 557592 526804
rect 547880 523728 547932 523734
rect 547880 523670 547932 523676
rect 543004 523116 543056 523122
rect 543004 523058 543056 523064
rect 542360 509244 542412 509250
rect 542360 509186 542412 509192
rect 542372 503674 542400 509186
rect 542360 503668 542412 503674
rect 542360 503610 542412 503616
rect 543016 500954 543044 523058
rect 545764 522300 545816 522306
rect 545764 522242 545816 522248
rect 545776 512281 545804 522242
rect 547892 521778 547920 523670
rect 557540 523116 557592 523122
rect 557540 523058 557592 523064
rect 557552 521778 557580 523058
rect 567200 523048 567252 523054
rect 567200 522990 567252 522996
rect 567212 521778 567240 522990
rect 547892 521750 548044 521778
rect 557552 521750 557704 521778
rect 567212 521750 567364 521778
rect 545762 512272 545818 512281
rect 545762 512207 545818 512216
rect 547892 502030 548044 502058
rect 557552 502030 557704 502058
rect 567212 502030 567364 502058
rect 543004 500948 543056 500954
rect 543004 500890 543056 500896
rect 547892 500818 547920 502030
rect 547880 500812 547932 500818
rect 547880 500754 547932 500760
rect 557552 500682 557580 502030
rect 567212 500886 567240 502030
rect 567200 500880 567252 500886
rect 567200 500822 567252 500828
rect 557540 500676 557592 500682
rect 557540 500618 557592 500624
rect 547880 497480 547932 497486
rect 547880 497422 547932 497428
rect 543004 496936 543056 496942
rect 543004 496878 543056 496884
rect 542358 484664 542414 484673
rect 542358 484599 542414 484608
rect 542372 476066 542400 484599
rect 542360 476060 542412 476066
rect 542360 476002 542412 476008
rect 543016 475930 543044 496878
rect 547892 494850 547920 497422
rect 557540 496936 557592 496942
rect 557540 496878 557592 496884
rect 557552 494850 557580 496878
rect 567200 496868 567252 496874
rect 567200 496810 567252 496816
rect 567212 494850 567240 496810
rect 547892 494822 548044 494850
rect 557552 494822 557704 494850
rect 567212 494822 567364 494850
rect 545764 494760 545816 494766
rect 545764 494702 545816 494708
rect 545776 485353 545804 494702
rect 545762 485344 545818 485353
rect 545762 485279 545818 485288
rect 543004 475924 543056 475930
rect 543004 475866 543056 475872
rect 547892 475102 548044 475130
rect 557552 475102 557704 475130
rect 567212 475102 567364 475130
rect 547892 473210 547920 475102
rect 547880 473204 547932 473210
rect 547880 473146 547932 473152
rect 557552 473074 557580 475102
rect 567212 473278 567240 475102
rect 567200 473272 567252 473278
rect 567200 473214 567252 473220
rect 557540 473068 557592 473074
rect 557540 473010 557592 473016
rect 547880 469872 547932 469878
rect 547880 469814 547932 469820
rect 543004 469328 543056 469334
rect 543004 469270 543056 469276
rect 542360 466472 542412 466478
rect 542360 466414 542412 466420
rect 542372 457609 542400 466414
rect 542358 457600 542414 457609
rect 542358 457535 542414 457544
rect 543016 448526 543044 469270
rect 545764 468512 545816 468518
rect 545764 468454 545816 468460
rect 545776 458289 545804 468454
rect 547892 467786 547920 469814
rect 557540 469328 557592 469334
rect 557540 469270 557592 469276
rect 557552 467786 557580 469270
rect 567200 469260 567252 469266
rect 567200 469202 567252 469208
rect 567212 467786 567240 469202
rect 547892 467758 548044 467786
rect 557552 467758 557704 467786
rect 567212 467758 567364 467786
rect 545762 458280 545818 458289
rect 545762 458215 545818 458224
rect 543004 448520 543056 448526
rect 543004 448462 543056 448468
rect 547892 448038 548044 448066
rect 557552 448038 557704 448066
rect 567212 448038 567364 448066
rect 547892 445602 547920 448038
rect 547880 445596 547932 445602
rect 547880 445538 547932 445544
rect 557552 445466 557580 448038
rect 567212 445670 567240 448038
rect 567200 445664 567252 445670
rect 567200 445606 567252 445612
rect 557540 445460 557592 445466
rect 557540 445402 557592 445408
rect 547880 443692 547932 443698
rect 547880 443634 547932 443640
rect 543004 443080 543056 443086
rect 543004 443022 543056 443028
rect 542360 440292 542412 440298
rect 542360 440234 542412 440240
rect 542372 430681 542400 440234
rect 542358 430672 542414 430681
rect 542358 430607 542414 430616
rect 543016 421734 543044 443022
rect 547892 440994 547920 443634
rect 557540 443080 557592 443086
rect 557540 443022 557592 443028
rect 557552 440994 557580 443022
rect 567200 443012 567252 443018
rect 567200 442954 567252 442960
rect 567212 440994 567240 442954
rect 547892 440966 548044 440994
rect 557552 440966 557704 440994
rect 567212 440966 567364 440994
rect 545764 440904 545816 440910
rect 545764 440846 545816 440852
rect 545776 431905 545804 440846
rect 545762 431896 545818 431905
rect 545762 431831 545818 431840
rect 543004 421728 543056 421734
rect 543004 421670 543056 421676
rect 547892 421110 548044 421138
rect 557552 421110 557704 421138
rect 567212 421110 567364 421138
rect 547892 419354 547920 421110
rect 547880 419348 547932 419354
rect 547880 419290 547932 419296
rect 557552 419218 557580 421110
rect 567212 419422 567240 421110
rect 567200 419416 567252 419422
rect 567200 419358 567252 419364
rect 557540 419212 557592 419218
rect 557540 419154 557592 419160
rect 547880 416084 547932 416090
rect 547880 416026 547932 416032
rect 543004 415540 543056 415546
rect 543004 415482 543056 415488
rect 542358 403608 542414 403617
rect 542358 403543 542414 403552
rect 542372 394670 542400 403543
rect 542360 394664 542412 394670
rect 542360 394606 542412 394612
rect 543016 391950 543044 415482
rect 545764 414724 545816 414730
rect 545764 414666 545816 414672
rect 545776 404297 545804 414666
rect 547892 413794 547920 416026
rect 557540 415540 557592 415546
rect 557540 415482 557592 415488
rect 557552 413794 557580 415482
rect 567200 415472 567252 415478
rect 567200 415414 567252 415420
rect 567212 413794 567240 415414
rect 547892 413766 548044 413794
rect 557552 413766 557704 413794
rect 567212 413766 567364 413794
rect 545762 404288 545818 404297
rect 545762 404223 545818 404232
rect 547892 394046 548044 394074
rect 557552 394046 557704 394074
rect 567212 394046 567364 394074
rect 543004 391944 543056 391950
rect 543004 391886 543056 391892
rect 547892 391814 547920 394046
rect 547880 391808 547932 391814
rect 547880 391750 547932 391756
rect 557552 391678 557580 394046
rect 567212 391882 567240 394046
rect 567200 391876 567252 391882
rect 567200 391818 567252 391824
rect 557540 391672 557592 391678
rect 557540 391614 557592 391620
rect 547880 389836 547932 389842
rect 547880 389778 547932 389784
rect 543004 389292 543056 389298
rect 543004 389234 543056 389240
rect 543016 365702 543044 389234
rect 545764 387116 545816 387122
rect 545764 387058 545816 387064
rect 545776 377913 545804 387058
rect 547892 386730 547920 389778
rect 557540 389292 557592 389298
rect 557540 389234 557592 389240
rect 557552 386730 557580 389234
rect 567200 389224 567252 389230
rect 567200 389166 567252 389172
rect 567212 386730 567240 389166
rect 547892 386702 548044 386730
rect 557552 386702 557704 386730
rect 567212 386702 567364 386730
rect 545762 377904 545818 377913
rect 545762 377839 545818 377848
rect 547892 367118 548044 367146
rect 557552 367118 557704 367146
rect 567212 367118 567364 367146
rect 543004 365696 543056 365702
rect 543004 365638 543056 365644
rect 547892 365566 547920 367118
rect 547880 365560 547932 365566
rect 547880 365502 547932 365508
rect 557552 365430 557580 367118
rect 567212 365634 567240 367118
rect 567200 365628 567252 365634
rect 567200 365570 567252 365576
rect 557540 365424 557592 365430
rect 557540 365366 557592 365372
rect 547880 362228 547932 362234
rect 547880 362170 547932 362176
rect 543004 361684 543056 361690
rect 543004 361626 543056 361632
rect 542358 349616 542414 349625
rect 542358 349551 542414 349560
rect 542372 340882 542400 349551
rect 542360 340876 542412 340882
rect 542360 340818 542412 340824
rect 543016 340746 543044 361626
rect 547892 359802 547920 362170
rect 557540 361684 557592 361690
rect 557540 361626 557592 361632
rect 557552 359802 557580 361626
rect 567200 361616 567252 361622
rect 567200 361558 567252 361564
rect 567212 359802 567240 361558
rect 547892 359774 548044 359802
rect 557552 359774 557704 359802
rect 567212 359774 567364 359802
rect 545764 359508 545816 359514
rect 545764 359450 545816 359456
rect 545776 350305 545804 359450
rect 545762 350296 545818 350305
rect 545762 350231 545818 350240
rect 543004 340740 543056 340746
rect 543004 340682 543056 340688
rect 547892 340054 548044 340082
rect 557552 340054 557704 340082
rect 567212 340054 567364 340082
rect 547892 337958 547920 340054
rect 547880 337952 547932 337958
rect 547880 337894 547932 337900
rect 557552 337822 557580 340054
rect 567212 338026 567240 340054
rect 567200 338020 567252 338026
rect 567200 337962 567252 337968
rect 557540 337816 557592 337822
rect 557540 337758 557592 337764
rect 547880 336048 547932 336054
rect 547880 335990 547932 335996
rect 543004 335436 543056 335442
rect 543004 335378 543056 335384
rect 542358 322008 542414 322017
rect 542358 321943 542414 321952
rect 542372 314634 542400 321943
rect 542360 314628 542412 314634
rect 542360 314570 542412 314576
rect 543016 311846 543044 335378
rect 545764 333260 545816 333266
rect 545764 333202 545816 333208
rect 545776 323921 545804 333202
rect 547892 332874 547920 335990
rect 557540 335436 557592 335442
rect 557540 335378 557592 335384
rect 557552 332874 557580 335378
rect 567200 335368 567252 335374
rect 567200 335310 567252 335316
rect 567212 332874 567240 335310
rect 547892 332846 548044 332874
rect 557552 332846 557704 332874
rect 567212 332846 567364 332874
rect 545762 323912 545818 323921
rect 545762 323847 545818 323856
rect 547892 313126 548044 313154
rect 557552 313126 557704 313154
rect 567212 313126 567364 313154
rect 543004 311840 543056 311846
rect 543004 311782 543056 311788
rect 547892 311710 547920 313126
rect 547880 311704 547932 311710
rect 547880 311646 547932 311652
rect 557552 311574 557580 313126
rect 567212 311778 567240 313126
rect 567200 311772 567252 311778
rect 567200 311714 567252 311720
rect 557540 311568 557592 311574
rect 557540 311510 557592 311516
rect 547880 308440 547932 308446
rect 547880 308382 547932 308388
rect 543004 307896 543056 307902
rect 543004 307838 543056 307844
rect 542358 295624 542414 295633
rect 542358 295559 542414 295568
rect 542372 287026 542400 295559
rect 542360 287020 542412 287026
rect 542360 286962 542412 286968
rect 543016 286822 543044 307838
rect 547892 305946 547920 308382
rect 557540 307896 557592 307902
rect 557540 307838 557592 307844
rect 557552 305946 557580 307838
rect 567200 307828 567252 307834
rect 567200 307770 567252 307776
rect 567212 305946 567240 307770
rect 547892 305918 548044 305946
rect 557552 305918 557704 305946
rect 567212 305918 567364 305946
rect 545764 305652 545816 305658
rect 545764 305594 545816 305600
rect 545776 296313 545804 305594
rect 545762 296304 545818 296313
rect 545762 296239 545818 296248
rect 543004 286816 543056 286822
rect 543004 286758 543056 286764
rect 547892 286062 548044 286090
rect 557552 286062 557704 286090
rect 567212 286062 567364 286090
rect 547892 284170 547920 286062
rect 547880 284164 547932 284170
rect 547880 284106 547932 284112
rect 557552 284034 557580 286062
rect 567212 284238 567240 286062
rect 567200 284232 567252 284238
rect 567200 284174 567252 284180
rect 557540 284028 557592 284034
rect 557540 283970 557592 283976
rect 547880 280832 547932 280838
rect 547880 280774 547932 280780
rect 543004 280288 543056 280294
rect 543004 280230 543056 280236
rect 542360 277432 542412 277438
rect 542360 277374 542412 277380
rect 542372 268569 542400 277374
rect 542358 268560 542414 268569
rect 542358 268495 542414 268504
rect 543016 256698 543044 280230
rect 545764 279472 545816 279478
rect 545764 279414 545816 279420
rect 545776 269793 545804 279414
rect 547892 278746 547920 280774
rect 557540 280288 557592 280294
rect 557540 280230 557592 280236
rect 557552 278746 557580 280230
rect 567200 280220 567252 280226
rect 567200 280162 567252 280168
rect 567212 278746 567240 280162
rect 547892 278718 548044 278746
rect 557552 278718 557704 278746
rect 567212 278718 567364 278746
rect 545762 269784 545818 269793
rect 545762 269719 545818 269728
rect 547892 259134 548044 259162
rect 557552 259134 557704 259162
rect 567212 259134 567364 259162
rect 543004 256692 543056 256698
rect 543004 256634 543056 256640
rect 547892 256562 547920 259134
rect 547880 256556 547932 256562
rect 547880 256498 547932 256504
rect 557552 256426 557580 259134
rect 567212 256630 567240 259134
rect 567200 256624 567252 256630
rect 567200 256566 567252 256572
rect 557540 256420 557592 256426
rect 557540 256362 557592 256368
rect 547880 254584 547932 254590
rect 547880 254526 547932 254532
rect 543004 254040 543056 254046
rect 543004 253982 543056 253988
rect 542360 251252 542412 251258
rect 542360 251194 542412 251200
rect 542372 241641 542400 251194
rect 542358 241632 542414 241641
rect 542358 241567 542414 241576
rect 543016 233170 543044 253982
rect 545764 251864 545816 251870
rect 545764 251806 545816 251812
rect 547892 251818 547920 254526
rect 557540 254040 557592 254046
rect 557540 253982 557592 253988
rect 557552 251818 557580 253982
rect 567200 253972 567252 253978
rect 567200 253914 567252 253920
rect 567212 251818 567240 253914
rect 545776 242321 545804 251806
rect 547892 251790 548044 251818
rect 557552 251790 557704 251818
rect 567212 251790 567364 251818
rect 545762 242312 545818 242321
rect 545762 242247 545818 242256
rect 543004 233164 543056 233170
rect 543004 233106 543056 233112
rect 547892 232070 548044 232098
rect 557552 232070 557704 232098
rect 567212 232070 567364 232098
rect 547892 230314 547920 232070
rect 547880 230308 547932 230314
rect 547880 230250 547932 230256
rect 557552 230178 557580 232070
rect 567212 230382 567240 232070
rect 567200 230376 567252 230382
rect 567200 230318 567252 230324
rect 557540 230172 557592 230178
rect 557540 230114 557592 230120
rect 547880 227044 547932 227050
rect 547880 226986 547932 226992
rect 543004 226432 543056 226438
rect 543004 226374 543056 226380
rect 542358 214568 542414 214577
rect 542358 214503 542414 214512
rect 542372 205630 542400 214503
rect 542360 205624 542412 205630
rect 542360 205566 542412 205572
rect 543016 205494 543044 226374
rect 545764 225616 545816 225622
rect 545764 225558 545816 225564
rect 545776 215257 545804 225558
rect 547892 224754 547920 226986
rect 557540 226432 557592 226438
rect 557540 226374 557592 226380
rect 557552 224754 557580 226374
rect 567200 226364 567252 226370
rect 567200 226306 567252 226312
rect 567212 224754 567240 226306
rect 547892 224726 548044 224754
rect 557552 224726 557704 224754
rect 567212 224726 567364 224754
rect 545762 215248 545818 215257
rect 545762 215183 545818 215192
rect 543004 205488 543056 205494
rect 543004 205430 543056 205436
rect 547892 205006 548044 205034
rect 557552 205006 557704 205034
rect 567212 205006 567364 205034
rect 547892 202706 547920 205006
rect 547880 202700 547932 202706
rect 547880 202642 547932 202648
rect 557552 202570 557580 205006
rect 567212 202774 567240 205006
rect 567200 202768 567252 202774
rect 567200 202710 567252 202716
rect 557540 202564 557592 202570
rect 557540 202506 557592 202512
rect 547880 200796 547932 200802
rect 547880 200738 547932 200744
rect 543004 200252 543056 200258
rect 543004 200194 543056 200200
rect 542358 187640 542414 187649
rect 542358 187575 542414 187584
rect 542372 179382 542400 187575
rect 542360 179376 542412 179382
rect 542360 179318 542412 179324
rect 543016 176662 543044 200194
rect 545764 198008 545816 198014
rect 545764 197950 545816 197956
rect 547892 197962 547920 200738
rect 557540 200252 557592 200258
rect 557540 200194 557592 200200
rect 557552 197962 557580 200194
rect 567200 200184 567252 200190
rect 567200 200126 567252 200132
rect 567212 197962 567240 200126
rect 545776 188329 545804 197950
rect 547892 197934 548044 197962
rect 557552 197934 557704 197962
rect 567212 197934 567364 197962
rect 545762 188320 545818 188329
rect 545762 188255 545818 188264
rect 547892 178078 548044 178106
rect 557552 178078 557704 178106
rect 567212 178078 567364 178106
rect 543004 176656 543056 176662
rect 543004 176598 543056 176604
rect 547892 176526 547920 178078
rect 547880 176520 547932 176526
rect 547880 176462 547932 176468
rect 557552 176390 557580 178078
rect 567212 176594 567240 178078
rect 567200 176588 567252 176594
rect 567200 176530 567252 176536
rect 557540 176384 557592 176390
rect 557540 176326 557592 176332
rect 547880 173188 547932 173194
rect 547880 173130 547932 173136
rect 543004 172644 543056 172650
rect 543004 172586 543056 172592
rect 542358 160576 542414 160585
rect 542358 160511 542414 160520
rect 542372 151774 542400 160511
rect 542360 151768 542412 151774
rect 542360 151710 542412 151716
rect 543016 151638 543044 172586
rect 547892 170898 547920 173130
rect 557540 172644 557592 172650
rect 557540 172586 557592 172592
rect 557552 170898 557580 172586
rect 567200 172576 567252 172582
rect 567200 172518 567252 172524
rect 567212 170898 567240 172518
rect 547892 170870 548044 170898
rect 557552 170870 557704 170898
rect 567212 170870 567364 170898
rect 545764 170400 545816 170406
rect 545764 170342 545816 170348
rect 545776 161265 545804 170342
rect 545762 161256 545818 161265
rect 545762 161191 545818 161200
rect 543004 151632 543056 151638
rect 543004 151574 543056 151580
rect 547892 151014 548044 151042
rect 557552 151014 557704 151042
rect 567212 151014 567364 151042
rect 547892 148918 547920 151014
rect 547880 148912 547932 148918
rect 547880 148854 547932 148860
rect 557552 148782 557580 151014
rect 567212 148986 567240 151014
rect 567200 148980 567252 148986
rect 567200 148922 567252 148928
rect 557540 148776 557592 148782
rect 557540 148718 557592 148724
rect 547880 146940 547932 146946
rect 547880 146882 547932 146888
rect 543004 146396 543056 146402
rect 543004 146338 543056 146344
rect 542358 133648 542414 133657
rect 542358 133583 542414 133592
rect 542372 125594 542400 133583
rect 542360 125588 542412 125594
rect 542360 125530 542412 125536
rect 543016 122806 543044 146338
rect 545764 144220 545816 144226
rect 545764 144162 545816 144168
rect 545776 134337 545804 144162
rect 547892 143834 547920 146882
rect 557540 146396 557592 146402
rect 557540 146338 557592 146344
rect 557552 143834 557580 146338
rect 567200 146328 567252 146334
rect 567200 146270 567252 146276
rect 567212 143834 567240 146270
rect 547892 143806 548044 143834
rect 557552 143806 557704 143834
rect 567212 143806 567364 143834
rect 545762 134328 545818 134337
rect 545762 134263 545818 134272
rect 547892 124086 548044 124114
rect 557552 124086 557704 124114
rect 567212 124086 567364 124114
rect 543004 122800 543056 122806
rect 543004 122742 543056 122748
rect 547892 122670 547920 124086
rect 557552 122738 557580 124086
rect 557540 122732 557592 122738
rect 557540 122674 557592 122680
rect 547880 122664 547932 122670
rect 547880 122606 547932 122612
rect 567212 122534 567240 124086
rect 567200 122528 567252 122534
rect 567200 122470 567252 122476
rect 547880 119400 547932 119406
rect 547880 119342 547932 119348
rect 543004 118788 543056 118794
rect 543004 118730 543056 118736
rect 542358 106584 542414 106593
rect 542358 106519 542414 106528
rect 542372 97986 542400 106519
rect 542360 97980 542412 97986
rect 542360 97922 542412 97928
rect 543016 97850 543044 118730
rect 547892 116770 547920 119342
rect 557540 118788 557592 118794
rect 557540 118730 557592 118736
rect 557552 116770 557580 118730
rect 567200 118720 567252 118726
rect 567200 118662 567252 118668
rect 567212 116770 567240 118662
rect 547892 116742 548044 116770
rect 557552 116742 557704 116770
rect 567212 116742 567364 116770
rect 545764 116612 545816 116618
rect 545764 116554 545816 116560
rect 545776 107273 545804 116554
rect 545762 107264 545818 107273
rect 545762 107199 545818 107208
rect 543004 97844 543056 97850
rect 543004 97786 543056 97792
rect 547892 97022 548044 97050
rect 557552 97022 557704 97050
rect 567212 97022 567364 97050
rect 547892 95062 547920 97022
rect 547880 95056 547932 95062
rect 547880 94998 547932 95004
rect 557552 94926 557580 97022
rect 567212 95130 567240 97022
rect 567200 95124 567252 95130
rect 567200 95066 567252 95072
rect 557540 94920 557592 94926
rect 557540 94862 557592 94868
rect 547880 91792 547932 91798
rect 547880 91734 547932 91740
rect 543004 91180 543056 91186
rect 543004 91122 543056 91128
rect 542358 79656 542414 79665
rect 542358 79591 542414 79600
rect 542372 71738 542400 79591
rect 542360 71732 542412 71738
rect 542360 71674 542412 71680
rect 543016 69018 543044 91122
rect 545764 90364 545816 90370
rect 545764 90306 545816 90312
rect 545776 80345 545804 90306
rect 547892 89842 547920 91734
rect 557540 91180 557592 91186
rect 557540 91122 557592 91128
rect 557552 89842 557580 91122
rect 567200 91112 567252 91118
rect 567200 91054 567252 91060
rect 567212 89842 567240 91054
rect 547892 89814 548044 89842
rect 557552 89814 557704 89842
rect 567212 89814 567364 89842
rect 545762 80336 545818 80345
rect 545762 80271 545818 80280
rect 547892 70094 548044 70122
rect 557552 70094 557704 70122
rect 567212 70094 567364 70122
rect 543004 69012 543056 69018
rect 543004 68954 543056 68960
rect 547892 68882 547920 70094
rect 547880 68876 547932 68882
rect 547880 68818 547932 68824
rect 557552 68746 557580 70094
rect 567212 68950 567240 70094
rect 567200 68944 567252 68950
rect 567200 68886 567252 68892
rect 557540 68740 557592 68746
rect 557540 68682 557592 68688
rect 547880 65544 547932 65550
rect 547880 65486 547932 65492
rect 543004 65000 543056 65006
rect 543004 64942 543056 64948
rect 542360 62144 542412 62150
rect 542360 62086 542412 62092
rect 542372 52601 542400 62086
rect 542358 52592 542414 52601
rect 542358 52527 542414 52536
rect 543016 44062 543044 64942
rect 547892 62914 547920 65486
rect 557540 65000 557592 65006
rect 557540 64942 557592 64948
rect 557552 62914 557580 64942
rect 567200 64932 567252 64938
rect 567200 64874 567252 64880
rect 567212 62914 567240 64874
rect 547892 62886 548044 62914
rect 557552 62886 557704 62914
rect 567212 62886 567364 62914
rect 545764 62824 545816 62830
rect 545764 62766 545816 62772
rect 545776 53281 545804 62766
rect 545762 53272 545818 53281
rect 545762 53207 545818 53216
rect 543004 44056 543056 44062
rect 543004 43998 543056 44004
rect 547892 43030 548044 43058
rect 557552 43030 557704 43058
rect 567212 43030 567364 43058
rect 547892 41274 547920 43030
rect 547880 41268 547932 41274
rect 547880 41210 547932 41216
rect 557552 41138 557580 43030
rect 567212 41342 567240 43030
rect 567200 41336 567252 41342
rect 567200 41278 567252 41284
rect 557540 41132 557592 41138
rect 557540 41074 557592 41080
rect 567856 38010 567884 670686
rect 569972 665174 570000 673503
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 569960 665168 570012 665174
rect 569960 665110 570012 665116
rect 569960 655648 570012 655654
rect 569960 655590 570012 655596
rect 569972 646649 570000 655590
rect 569958 646640 570014 646649
rect 569958 646575 570014 646584
rect 569958 619576 570014 619585
rect 569958 619511 570014 619520
rect 567936 616888 567988 616894
rect 567936 616830 567988 616836
rect 567844 38004 567896 38010
rect 567844 37946 567896 37952
rect 547972 37936 548024 37942
rect 547972 37878 548024 37884
rect 543004 37392 543056 37398
rect 543004 37334 543056 37340
rect 542360 34536 542412 34542
rect 542360 34478 542412 34484
rect 542372 25673 542400 34478
rect 542358 25664 542414 25673
rect 542358 25599 542414 25608
rect 543016 16590 543044 37334
rect 547144 37324 547196 37330
rect 547144 37266 547196 37272
rect 545764 36644 545816 36650
rect 545764 36586 545816 36592
rect 545776 26353 545804 36586
rect 545762 26344 545818 26353
rect 545762 26279 545818 26288
rect 543004 16584 543056 16590
rect 543004 16526 543056 16532
rect 547156 13462 547184 37266
rect 547984 36122 548012 37878
rect 557540 37392 557592 37398
rect 557540 37334 557592 37340
rect 547984 36094 548058 36122
rect 548030 35972 548058 36094
rect 557552 35986 557580 37334
rect 567200 37324 567252 37330
rect 567200 37266 567252 37272
rect 557552 35958 557704 35986
rect 567212 35894 567240 37266
rect 567350 35894 567378 35972
rect 567212 35866 567378 35894
rect 547892 16102 548044 16130
rect 557552 16102 557704 16130
rect 567212 16102 567364 16130
rect 547892 13598 547920 16102
rect 557552 13666 557580 16102
rect 557540 13660 557592 13666
rect 557540 13602 557592 13608
rect 547880 13592 547932 13598
rect 547880 13534 547932 13540
rect 567212 13530 567240 16102
rect 567200 13524 567252 13530
rect 567200 13466 567252 13472
rect 547144 13456 547196 13462
rect 547144 13398 547196 13404
rect 567948 13394 567976 616830
rect 569972 611250 570000 619511
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 569960 611244 570012 611250
rect 569960 611186 570012 611192
rect 569958 592648 570014 592657
rect 569958 592583 570014 592592
rect 569972 583642 570000 592583
rect 569960 583636 570012 583642
rect 569960 583578 570012 583584
rect 569958 565584 570014 565593
rect 569958 565519 570014 565528
rect 569972 557462 570000 565519
rect 580262 564360 580318 564369
rect 580262 564295 580318 564304
rect 569960 557456 570012 557462
rect 569960 557398 570012 557404
rect 569958 538656 570014 538665
rect 569958 538591 570014 538600
rect 569972 529854 570000 538591
rect 569960 529848 570012 529854
rect 569960 529790 570012 529796
rect 569960 520328 570012 520334
rect 569960 520270 570012 520276
rect 569972 511601 570000 520270
rect 569958 511592 570014 511601
rect 569958 511527 570014 511536
rect 569958 484664 570014 484673
rect 569958 484599 570014 484608
rect 569972 475998 570000 484599
rect 569960 475992 570012 475998
rect 569960 475934 570012 475940
rect 569960 466540 570012 466546
rect 569960 466482 570012 466488
rect 569972 457609 570000 466482
rect 569958 457600 570014 457609
rect 569958 457535 570014 457544
rect 569958 430672 570014 430681
rect 569958 430607 570014 430616
rect 569972 422278 570000 430607
rect 569960 422272 570012 422278
rect 569960 422214 570012 422220
rect 569958 403608 570014 403617
rect 569958 403543 570014 403552
rect 569972 394602 570000 403543
rect 569960 394596 570012 394602
rect 569960 394538 570012 394544
rect 569958 376000 570014 376009
rect 569958 375935 570014 375944
rect 569972 368422 570000 375935
rect 569960 368416 570012 368422
rect 569960 368358 570012 368364
rect 569958 349616 570014 349625
rect 569958 349551 570014 349560
rect 569972 340814 570000 349551
rect 569960 340808 570012 340814
rect 569960 340750 570012 340756
rect 569958 322008 570014 322017
rect 569958 321943 570014 321952
rect 569972 314566 570000 321943
rect 569960 314560 570012 314566
rect 569960 314502 570012 314508
rect 569958 295624 570014 295633
rect 569958 295559 570014 295568
rect 569972 286958 570000 295559
rect 569960 286952 570012 286958
rect 569960 286894 570012 286900
rect 569960 277500 570012 277506
rect 569960 277442 570012 277448
rect 569972 268569 570000 277442
rect 569958 268560 570014 268569
rect 569958 268495 570014 268504
rect 569958 241632 570014 241641
rect 569958 241567 570014 241576
rect 569972 233238 570000 241567
rect 569960 233232 570012 233238
rect 569960 233174 570012 233180
rect 569958 214568 570014 214577
rect 569958 214503 570014 214512
rect 569972 205562 570000 214503
rect 569960 205556 570012 205562
rect 569960 205498 570012 205504
rect 569958 187640 570014 187649
rect 569958 187575 570014 187584
rect 569972 179314 570000 187575
rect 569960 179308 570012 179314
rect 569960 179250 570012 179256
rect 569958 160576 570014 160585
rect 569958 160511 570014 160520
rect 569972 151706 570000 160511
rect 569960 151700 570012 151706
rect 569960 151642 570012 151648
rect 569958 133648 570014 133657
rect 569958 133583 570014 133592
rect 569972 125526 570000 133583
rect 569960 125520 570012 125526
rect 569960 125462 570012 125468
rect 569958 106584 570014 106593
rect 569958 106519 570014 106528
rect 569972 97918 570000 106519
rect 569960 97912 570012 97918
rect 569960 97854 570012 97860
rect 569960 88392 570012 88398
rect 569960 88334 570012 88340
rect 569972 79665 570000 88334
rect 569958 79656 570014 79665
rect 569958 79591 570014 79600
rect 569958 52592 570014 52601
rect 569958 52527 570014 52536
rect 569972 44130 570000 52527
rect 569960 44124 570012 44130
rect 569960 44066 570012 44072
rect 580276 36582 580304 564295
rect 580264 36576 580316 36582
rect 580264 36518 580316 36524
rect 569960 34604 570012 34610
rect 569960 34546 570012 34552
rect 569972 25673 570000 34546
rect 569958 25664 570014 25673
rect 569958 25599 570014 25608
rect 567936 13388 567988 13394
rect 567936 13330 567988 13336
rect 541624 13320 541676 13326
rect 541624 13262 541676 13268
rect 3424 13116 3476 13122
rect 3424 13058 3476 13064
rect 43720 13116 43772 13122
rect 43720 13058 43772 13064
rect 3436 6497 3464 13058
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3146 632068 3148 632088
rect 3148 632068 3200 632088
rect 3200 632068 3202 632088
rect 3146 632032 3202 632068
rect 3238 579944 3294 580000
rect 3422 527856 3478 527912
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 358400 3386 358456
rect 3054 306176 3110 306232
rect 3330 254108 3386 254144
rect 3330 254088 3332 254108
rect 3332 254088 3384 254108
rect 3384 254088 3386 254108
rect 3054 241032 3110 241088
rect 2962 188808 3018 188864
rect 3146 84632 3202 84688
rect 3330 58520 3386 58576
rect 3238 45464 3294 45520
rect 3514 475632 3570 475688
rect 3606 345344 3662 345400
rect 3698 293120 3754 293176
rect 3790 201864 3846 201920
rect 3422 19352 3478 19408
rect 3882 149776 3938 149832
rect 3974 136720 4030 136776
rect 4066 97552 4122 97608
rect 13726 674192 13782 674248
rect 13726 647264 13782 647320
rect 13726 620200 13782 620256
rect 13726 593272 13782 593328
rect 13726 566208 13782 566264
rect 13726 539280 13782 539336
rect 13726 512216 13782 512272
rect 13726 485288 13782 485344
rect 13726 458224 13782 458280
rect 13726 431296 13782 431352
rect 13726 404232 13782 404288
rect 13726 376760 13782 376816
rect 13726 350240 13782 350296
rect 13726 322904 13782 322960
rect 13726 296248 13782 296304
rect 13726 269184 13782 269240
rect 13726 242256 13782 242312
rect 13726 215192 13782 215248
rect 13726 188264 13782 188320
rect 11702 35808 11758 35864
rect 12438 32408 12494 32464
rect 13726 161200 13782 161256
rect 13726 134272 13782 134328
rect 13726 107208 13782 107264
rect 13726 80280 13782 80336
rect 13726 53216 13782 53272
rect 13726 29008 13782 29064
rect 13726 25608 13782 25664
rect 13174 22208 13230 22264
rect 12438 18808 12494 18864
rect 37922 673512 37978 673568
rect 37922 646584 37978 646640
rect 37922 619520 37978 619576
rect 37922 592592 37978 592648
rect 37922 565528 37978 565584
rect 37922 538600 37978 538656
rect 37922 511536 37978 511592
rect 37922 484608 37978 484664
rect 37922 457544 37978 457600
rect 37922 430616 37978 430672
rect 37922 403552 37978 403608
rect 37922 375944 37978 376000
rect 37922 349560 37978 349616
rect 37922 321952 37978 322008
rect 37922 295568 37978 295624
rect 37922 268504 37978 268560
rect 37922 241576 37978 241632
rect 37922 214512 37978 214568
rect 37922 187584 37978 187640
rect 37922 160520 37978 160576
rect 37922 133592 37978 133648
rect 37922 106528 37978 106584
rect 37922 79600 37978 79656
rect 37922 52536 37978 52592
rect 42706 674192 42762 674248
rect 42706 647264 42762 647320
rect 42706 620200 42762 620256
rect 42706 593272 42762 593328
rect 42706 566208 42762 566264
rect 42706 539280 42762 539336
rect 42706 512216 42762 512272
rect 42706 485288 42762 485344
rect 42706 458224 42762 458280
rect 42706 431296 42762 431352
rect 42706 404232 42762 404288
rect 42706 376760 42762 376816
rect 42706 350240 42762 350296
rect 42706 322904 42762 322960
rect 42706 296248 42762 296304
rect 42706 269184 42762 269240
rect 42706 242256 42762 242312
rect 42706 215192 42762 215248
rect 42706 188264 42762 188320
rect 42706 161200 42762 161256
rect 42706 134272 42762 134328
rect 42706 107208 42762 107264
rect 42706 80280 42762 80336
rect 42706 53216 42762 53272
rect 61290 36100 61346 36136
rect 61290 36080 61292 36100
rect 61292 36080 61344 36100
rect 61344 36080 61346 36100
rect 63498 33088 63554 33144
rect 63590 29688 63646 29744
rect 63498 26288 63554 26344
rect 63498 19488 63554 19544
rect 64234 22888 64290 22944
rect 64418 16088 64474 16144
rect 66258 673512 66314 673568
rect 66258 646584 66314 646640
rect 66258 619520 66314 619576
rect 66258 592592 66314 592648
rect 66258 565528 66314 565584
rect 66258 538600 66314 538656
rect 66258 511536 66314 511592
rect 66258 484608 66314 484664
rect 66258 457544 66314 457600
rect 66258 430616 66314 430672
rect 66258 403552 66314 403608
rect 66258 375944 66314 376000
rect 66258 349560 66314 349616
rect 66258 321952 66314 322008
rect 66258 295568 66314 295624
rect 66258 268504 66314 268560
rect 66258 241576 66314 241632
rect 66258 214512 66314 214568
rect 66258 187584 66314 187640
rect 66258 160520 66314 160576
rect 66258 133592 66314 133648
rect 66258 106528 66314 106584
rect 66258 79600 66314 79656
rect 66258 52536 66314 52592
rect 70306 673784 70362 673840
rect 70306 647264 70362 647320
rect 93858 673512 93914 673568
rect 97906 674192 97962 674248
rect 126886 674192 126942 674248
rect 121458 673512 121514 673568
rect 154486 674192 154542 674248
rect 149058 673512 149114 673568
rect 178038 673512 178094 673568
rect 182086 674192 182142 674248
rect 209686 674192 209742 674248
rect 205638 674056 205694 674112
rect 233238 673512 233294 673568
rect 93858 646584 93914 646640
rect 97906 647264 97962 647320
rect 126886 647264 126942 647320
rect 121458 646584 121514 646640
rect 154486 647264 154542 647320
rect 149058 646584 149114 646640
rect 178038 646584 178094 646640
rect 182086 647264 182142 647320
rect 209686 647264 209742 647320
rect 205638 646584 205694 646640
rect 233238 646584 233294 646640
rect 70306 620200 70362 620256
rect 70306 593272 70362 593328
rect 93858 619520 93914 619576
rect 97906 620200 97962 620256
rect 126886 620200 126942 620256
rect 121458 619520 121514 619576
rect 154486 620200 154542 620256
rect 149058 619520 149114 619576
rect 178038 619520 178094 619576
rect 182086 620200 182142 620256
rect 209686 620200 209742 620256
rect 205638 619520 205694 619576
rect 233238 619520 233294 619576
rect 93858 592592 93914 592648
rect 97906 593272 97962 593328
rect 126886 593272 126942 593328
rect 121458 592592 121514 592648
rect 154486 593272 154542 593328
rect 149058 592592 149114 592648
rect 178038 592592 178094 592648
rect 182086 593272 182142 593328
rect 209686 593272 209742 593328
rect 205638 592592 205694 592648
rect 233238 592592 233294 592648
rect 70306 566208 70362 566264
rect 70306 539280 70362 539336
rect 93858 565528 93914 565584
rect 97906 566208 97962 566264
rect 126886 566208 126942 566264
rect 121458 565528 121514 565584
rect 154486 566208 154542 566264
rect 149058 565528 149114 565584
rect 178038 565528 178094 565584
rect 182086 566208 182142 566264
rect 209686 566208 209742 566264
rect 205638 565528 205694 565584
rect 233238 565528 233294 565584
rect 93858 538600 93914 538656
rect 97906 539280 97962 539336
rect 126886 539280 126942 539336
rect 121458 538600 121514 538656
rect 154486 539280 154542 539336
rect 149058 538600 149114 538656
rect 178038 538600 178094 538656
rect 182086 539280 182142 539336
rect 209686 539280 209742 539336
rect 205638 538600 205694 538656
rect 233238 538600 233294 538656
rect 70306 512216 70362 512272
rect 70306 484744 70362 484800
rect 93858 511536 93914 511592
rect 97906 512216 97962 512272
rect 126886 512216 126942 512272
rect 121458 511536 121514 511592
rect 154486 512216 154542 512272
rect 149058 511536 149114 511592
rect 178038 511536 178094 511592
rect 182086 512216 182142 512272
rect 209686 512216 209742 512272
rect 205638 511536 205694 511592
rect 233238 511536 233294 511592
rect 93858 484608 93914 484664
rect 97906 485288 97962 485344
rect 126886 485288 126942 485344
rect 121458 484608 121514 484664
rect 154486 485288 154542 485344
rect 149058 484608 149114 484664
rect 178038 484608 178094 484664
rect 182086 485288 182142 485344
rect 209686 485288 209742 485344
rect 205638 484472 205694 484528
rect 233238 484608 233294 484664
rect 70306 458224 70362 458280
rect 70306 430752 70362 430808
rect 93858 457544 93914 457600
rect 97906 458224 97962 458280
rect 126886 458224 126942 458280
rect 121458 457544 121514 457600
rect 154486 458224 154542 458280
rect 149058 457544 149114 457600
rect 178038 457544 178094 457600
rect 182086 458224 182142 458280
rect 209686 458224 209742 458280
rect 205638 457544 205694 457600
rect 233238 457544 233294 457600
rect 93858 430616 93914 430672
rect 97906 431296 97962 431352
rect 126886 431296 126942 431352
rect 121458 430616 121514 430672
rect 154486 431296 154542 431352
rect 149058 430616 149114 430672
rect 178038 430616 178094 430672
rect 182086 431296 182142 431352
rect 209686 431296 209742 431352
rect 205638 431160 205694 431216
rect 233238 430616 233294 430672
rect 70306 404232 70362 404288
rect 93858 403552 93914 403608
rect 97906 404232 97962 404288
rect 126886 404232 126942 404288
rect 121458 403552 121514 403608
rect 154486 404232 154542 404288
rect 149058 403552 149114 403608
rect 178038 403552 178094 403608
rect 182086 404232 182142 404288
rect 209686 404232 209742 404288
rect 205638 403552 205694 403608
rect 233238 403552 233294 403608
rect 70306 376760 70362 376816
rect 70306 350240 70362 350296
rect 93858 375944 93914 376000
rect 97906 376760 97962 376816
rect 126886 376760 126942 376816
rect 121458 375944 121514 376000
rect 154486 376760 154542 376816
rect 149058 375944 149114 376000
rect 178038 375944 178094 376000
rect 182086 376760 182142 376816
rect 209686 377032 209742 377088
rect 205638 375944 205694 376000
rect 233238 375944 233294 376000
rect 93858 349560 93914 349616
rect 97906 350240 97962 350296
rect 126886 350240 126942 350296
rect 121458 349560 121514 349616
rect 154486 350240 154542 350296
rect 149058 349560 149114 349616
rect 178038 349560 178094 349616
rect 182086 350240 182142 350296
rect 209686 350240 209742 350296
rect 205638 349560 205694 349616
rect 233238 349560 233294 349616
rect 70306 322904 70362 322960
rect 70306 296248 70362 296304
rect 93858 321952 93914 322008
rect 97906 322904 97962 322960
rect 126886 322904 126942 322960
rect 121458 321952 121514 322008
rect 154486 322904 154542 322960
rect 149058 321952 149114 322008
rect 178038 321952 178094 322008
rect 182086 322904 182142 322960
rect 209686 323856 209742 323912
rect 205638 321952 205694 322008
rect 233238 321952 233294 322008
rect 93858 295568 93914 295624
rect 97906 296248 97962 296304
rect 126886 296248 126942 296304
rect 121458 295568 121514 295624
rect 154486 296248 154542 296304
rect 149058 295568 149114 295624
rect 178038 295568 178094 295624
rect 182086 296248 182142 296304
rect 209686 296248 209742 296304
rect 205638 295568 205694 295624
rect 233238 295568 233294 295624
rect 70306 269728 70362 269784
rect 70306 242256 70362 242312
rect 93858 268504 93914 268560
rect 97906 269184 97962 269240
rect 126886 269184 126942 269240
rect 121458 268504 121514 268560
rect 154486 269184 154542 269240
rect 149058 268504 149114 268560
rect 178038 268504 178094 268560
rect 182086 269184 182142 269240
rect 209686 269184 209742 269240
rect 205638 269048 205694 269104
rect 233238 268504 233294 268560
rect 93858 241576 93914 241632
rect 97906 242256 97962 242312
rect 126886 242256 126942 242312
rect 121458 241576 121514 241632
rect 154486 242256 154542 242312
rect 149058 241576 149114 241632
rect 178038 241576 178094 241632
rect 182086 242256 182142 242312
rect 209686 242256 209742 242312
rect 205638 241576 205694 241632
rect 233238 241576 233294 241632
rect 70306 214648 70362 214704
rect 93858 214512 93914 214568
rect 97906 215192 97962 215248
rect 126886 215192 126942 215248
rect 121458 214512 121514 214568
rect 154486 215192 154542 215248
rect 149058 214512 149114 214568
rect 178038 214512 178094 214568
rect 182086 215192 182142 215248
rect 209686 215192 209742 215248
rect 205638 213968 205694 214024
rect 233238 214512 233294 214568
rect 70306 188264 70362 188320
rect 70306 161200 70362 161256
rect 93858 187584 93914 187640
rect 97906 188264 97962 188320
rect 126886 188264 126942 188320
rect 121458 187584 121514 187640
rect 154486 188264 154542 188320
rect 149058 187584 149114 187640
rect 178038 187584 178094 187640
rect 182086 188264 182142 188320
rect 209686 188264 209742 188320
rect 205638 187584 205694 187640
rect 233238 187584 233294 187640
rect 93858 160520 93914 160576
rect 97906 161200 97962 161256
rect 126886 161200 126942 161256
rect 121458 160520 121514 160576
rect 154486 161200 154542 161256
rect 149058 160520 149114 160576
rect 178038 160520 178094 160576
rect 182086 161200 182142 161256
rect 209686 161200 209742 161256
rect 205638 160520 205694 160576
rect 233238 160520 233294 160576
rect 70306 134272 70362 134328
rect 70306 107208 70362 107264
rect 93858 133592 93914 133648
rect 97906 134272 97962 134328
rect 126886 134272 126942 134328
rect 121458 133592 121514 133648
rect 154486 134272 154542 134328
rect 149058 133592 149114 133648
rect 178038 133592 178094 133648
rect 182086 134272 182142 134328
rect 209686 134272 209742 134328
rect 205638 133592 205694 133648
rect 233238 133592 233294 133648
rect 93858 106528 93914 106584
rect 97906 107208 97962 107264
rect 126886 107208 126942 107264
rect 121458 106528 121514 106584
rect 154486 107208 154542 107264
rect 149058 106528 149114 106584
rect 178038 106528 178094 106584
rect 182086 107208 182142 107264
rect 209686 107208 209742 107264
rect 205638 106528 205694 106584
rect 233238 106528 233294 106584
rect 70306 80280 70362 80336
rect 70306 53216 70362 53272
rect 93858 79600 93914 79656
rect 97906 80280 97962 80336
rect 126886 80280 126942 80336
rect 121458 79600 121514 79656
rect 154486 80280 154542 80336
rect 149058 79600 149114 79656
rect 178038 79600 178094 79656
rect 182086 80280 182142 80336
rect 209686 80280 209742 80336
rect 205638 79600 205694 79656
rect 233238 79600 233294 79656
rect 93858 52536 93914 52592
rect 97906 53216 97962 53272
rect 126886 53216 126942 53272
rect 121458 52536 121514 52592
rect 154486 53216 154542 53272
rect 149058 52536 149114 52592
rect 178038 52536 178094 52592
rect 182086 53216 182142 53272
rect 209686 53216 209742 53272
rect 205638 52536 205694 52592
rect 233238 52536 233294 52592
rect 238666 674192 238722 674248
rect 266266 674192 266322 674248
rect 262218 673512 262274 673568
rect 293866 674192 293922 674248
rect 289818 673512 289874 673568
rect 322846 674192 322902 674248
rect 317418 673512 317474 673568
rect 345018 673512 345074 673568
rect 350446 674192 350502 674248
rect 373998 673512 374054 673568
rect 378046 674192 378102 674248
rect 405646 674192 405702 674248
rect 401598 673512 401654 673568
rect 434626 674192 434682 674248
rect 429198 673512 429254 673568
rect 462226 674192 462282 674248
rect 458178 673512 458234 673568
rect 489826 674192 489882 674248
rect 485778 673512 485834 673568
rect 238666 647264 238722 647320
rect 266266 647264 266322 647320
rect 262218 646584 262274 646640
rect 293866 647264 293922 647320
rect 289818 646584 289874 646640
rect 322846 647264 322902 647320
rect 317418 646584 317474 646640
rect 345018 646584 345074 646640
rect 350446 647264 350502 647320
rect 373998 646584 374054 646640
rect 378046 647264 378102 647320
rect 405646 647264 405702 647320
rect 401598 646584 401654 646640
rect 434626 647264 434682 647320
rect 429198 646584 429254 646640
rect 462226 647264 462282 647320
rect 458178 646584 458234 646640
rect 489826 647264 489882 647320
rect 485778 646584 485834 646640
rect 238666 620200 238722 620256
rect 266266 620200 266322 620256
rect 262218 619520 262274 619576
rect 293866 620200 293922 620256
rect 289818 619520 289874 619576
rect 322846 620200 322902 620256
rect 317418 619520 317474 619576
rect 345018 619520 345074 619576
rect 350446 620200 350502 620256
rect 373998 619520 374054 619576
rect 378046 620200 378102 620256
rect 405646 620200 405702 620256
rect 401598 619520 401654 619576
rect 434626 620200 434682 620256
rect 429198 619520 429254 619576
rect 462226 620200 462282 620256
rect 458178 619520 458234 619576
rect 489826 620200 489882 620256
rect 485778 619520 485834 619576
rect 238666 593272 238722 593328
rect 238666 566208 238722 566264
rect 266266 593272 266322 593328
rect 262218 592592 262274 592648
rect 293866 593272 293922 593328
rect 289818 592592 289874 592648
rect 322846 593272 322902 593328
rect 317418 592592 317474 592648
rect 345018 592592 345074 592648
rect 350446 593272 350502 593328
rect 373998 592592 374054 592648
rect 378046 593272 378102 593328
rect 405646 593272 405702 593328
rect 401598 592592 401654 592648
rect 434626 593272 434682 593328
rect 429198 592592 429254 592648
rect 462226 593272 462282 593328
rect 458178 592592 458234 592648
rect 489826 593272 489882 593328
rect 485778 592592 485834 592648
rect 266266 566208 266322 566264
rect 262218 565528 262274 565584
rect 293866 566208 293922 566264
rect 289818 565528 289874 565584
rect 322846 566208 322902 566264
rect 317418 565528 317474 565584
rect 345018 565528 345074 565584
rect 350446 566208 350502 566264
rect 373998 565528 374054 565584
rect 378046 566208 378102 566264
rect 405646 566208 405702 566264
rect 401598 565528 401654 565584
rect 434626 566208 434682 566264
rect 429198 565528 429254 565584
rect 462226 566208 462282 566264
rect 458178 565528 458234 565584
rect 489826 566208 489882 566264
rect 485778 565528 485834 565584
rect 238666 539280 238722 539336
rect 238666 512216 238722 512272
rect 266266 539280 266322 539336
rect 262218 538600 262274 538656
rect 293866 539280 293922 539336
rect 289818 538600 289874 538656
rect 322846 539280 322902 539336
rect 317418 538600 317474 538656
rect 345018 538600 345074 538656
rect 350446 539280 350502 539336
rect 373998 538600 374054 538656
rect 378046 539280 378102 539336
rect 405646 539280 405702 539336
rect 401598 538600 401654 538656
rect 434626 539280 434682 539336
rect 429198 538600 429254 538656
rect 462226 539280 462282 539336
rect 458178 538600 458234 538656
rect 489826 539280 489882 539336
rect 485778 538600 485834 538656
rect 266266 512216 266322 512272
rect 262218 511536 262274 511592
rect 293866 512216 293922 512272
rect 289818 511536 289874 511592
rect 322846 512216 322902 512272
rect 317418 511536 317474 511592
rect 345018 511536 345074 511592
rect 350446 512216 350502 512272
rect 373998 511536 374054 511592
rect 378046 512216 378102 512272
rect 407854 512760 407910 512816
rect 401598 511536 401654 511592
rect 434626 512216 434682 512272
rect 429198 511536 429254 511592
rect 462226 512216 462282 512272
rect 458178 511536 458234 511592
rect 489826 512216 489882 512272
rect 485778 511536 485834 511592
rect 238666 485288 238722 485344
rect 238666 458224 238722 458280
rect 266266 485288 266322 485344
rect 262218 484608 262274 484664
rect 293866 485288 293922 485344
rect 289818 484608 289874 484664
rect 322846 485288 322902 485344
rect 317418 484608 317474 484664
rect 345018 484608 345074 484664
rect 350446 485288 350502 485344
rect 373998 484608 374054 484664
rect 378046 485288 378102 485344
rect 405646 485288 405702 485344
rect 401598 484608 401654 484664
rect 434626 485288 434682 485344
rect 429198 484608 429254 484664
rect 462226 485288 462282 485344
rect 458178 484608 458234 484664
rect 489826 485288 489882 485344
rect 485778 484608 485834 484664
rect 266266 458224 266322 458280
rect 262218 457544 262274 457600
rect 293866 458224 293922 458280
rect 289818 457544 289874 457600
rect 322846 458224 322902 458280
rect 317418 457544 317474 457600
rect 345018 457544 345074 457600
rect 350446 458224 350502 458280
rect 373998 457544 374054 457600
rect 378046 458224 378102 458280
rect 405646 458224 405702 458280
rect 401598 457544 401654 457600
rect 434626 458224 434682 458280
rect 429198 457544 429254 457600
rect 462226 458224 462282 458280
rect 458178 457544 458234 457600
rect 489826 458224 489882 458280
rect 485778 457544 485834 457600
rect 238666 431296 238722 431352
rect 266266 431296 266322 431352
rect 262218 430616 262274 430672
rect 293866 431296 293922 431352
rect 289818 430616 289874 430672
rect 322846 431296 322902 431352
rect 317418 430616 317474 430672
rect 345018 430616 345074 430672
rect 350446 431296 350502 431352
rect 373998 430752 374054 430808
rect 378046 431296 378102 431352
rect 405646 431296 405702 431352
rect 401598 430616 401654 430672
rect 434626 431296 434682 431352
rect 429198 430616 429254 430672
rect 462226 431296 462282 431352
rect 458178 430616 458234 430672
rect 489826 431296 489882 431352
rect 485778 430616 485834 430672
rect 238666 404232 238722 404288
rect 238666 377032 238722 377088
rect 260746 375944 260802 376000
rect 266266 404232 266322 404288
rect 262218 403552 262274 403608
rect 293866 404232 293922 404288
rect 289818 403552 289874 403608
rect 322846 404232 322902 404288
rect 317418 403552 317474 403608
rect 345018 403552 345074 403608
rect 350446 404232 350502 404288
rect 373998 403552 374054 403608
rect 378046 404232 378102 404288
rect 405646 404232 405702 404288
rect 401598 403552 401654 403608
rect 434626 404232 434682 404288
rect 429198 403552 429254 403608
rect 462226 404232 462282 404288
rect 458178 403552 458234 403608
rect 489826 404232 489882 404288
rect 485778 403552 485834 403608
rect 266266 377032 266322 377088
rect 293866 376760 293922 376816
rect 289818 375944 289874 376000
rect 322846 376760 322902 376816
rect 317418 375944 317474 376000
rect 345018 375944 345074 376000
rect 350446 376760 350502 376816
rect 373998 375944 374054 376000
rect 378046 376760 378102 376816
rect 405646 376760 405702 376816
rect 401598 375944 401654 376000
rect 434626 376760 434682 376816
rect 429198 375944 429254 376000
rect 462226 376760 462282 376816
rect 458178 375944 458234 376000
rect 489826 377032 489882 377088
rect 485778 375944 485834 376000
rect 238666 350240 238722 350296
rect 238666 322904 238722 322960
rect 266266 350240 266322 350296
rect 262218 349560 262274 349616
rect 293866 350240 293922 350296
rect 289818 349560 289874 349616
rect 322846 350240 322902 350296
rect 317418 349560 317474 349616
rect 345018 349560 345074 349616
rect 350446 350240 350502 350296
rect 373998 349560 374054 349616
rect 378046 350240 378102 350296
rect 405646 350240 405702 350296
rect 401598 349560 401654 349616
rect 434626 350240 434682 350296
rect 429198 349560 429254 349616
rect 462226 350240 462282 350296
rect 458178 349560 458234 349616
rect 489826 350240 489882 350296
rect 485778 349560 485834 349616
rect 266266 323856 266322 323912
rect 262218 322768 262274 322824
rect 293866 322904 293922 322960
rect 289818 321952 289874 322008
rect 322846 322904 322902 322960
rect 317418 322768 317474 322824
rect 345018 321952 345074 322008
rect 350446 322904 350502 322960
rect 373998 321952 374054 322008
rect 378046 322904 378102 322960
rect 405646 323856 405702 323912
rect 401598 321952 401654 322008
rect 434626 322904 434682 322960
rect 429198 321952 429254 322008
rect 462226 323856 462282 323912
rect 458178 322768 458234 322824
rect 489826 322904 489882 322960
rect 485778 321952 485834 322008
rect 238666 296248 238722 296304
rect 238666 269184 238722 269240
rect 266266 296248 266322 296304
rect 262218 295568 262274 295624
rect 293866 296248 293922 296304
rect 289818 295568 289874 295624
rect 322846 296248 322902 296304
rect 317418 295568 317474 295624
rect 345018 295568 345074 295624
rect 350446 296248 350502 296304
rect 373998 295568 374054 295624
rect 378046 296248 378102 296304
rect 405646 296248 405702 296304
rect 401598 295568 401654 295624
rect 434626 296248 434682 296304
rect 429198 295568 429254 295624
rect 462226 296248 462282 296304
rect 458178 295568 458234 295624
rect 489826 296248 489882 296304
rect 485778 295568 485834 295624
rect 266266 269184 266322 269240
rect 262218 268504 262274 268560
rect 293866 269184 293922 269240
rect 289818 268504 289874 268560
rect 322846 269184 322902 269240
rect 317418 268504 317474 268560
rect 345018 268504 345074 268560
rect 350446 269184 350502 269240
rect 373998 269048 374054 269104
rect 378046 269184 378102 269240
rect 405646 269184 405702 269240
rect 401598 268504 401654 268560
rect 434626 269184 434682 269240
rect 429198 268504 429254 268560
rect 462226 269184 462282 269240
rect 458178 268504 458234 268560
rect 489826 269184 489882 269240
rect 485778 268504 485834 268560
rect 238666 242256 238722 242312
rect 266266 242256 266322 242312
rect 262218 241576 262274 241632
rect 293866 242256 293922 242312
rect 289818 241576 289874 241632
rect 322846 242256 322902 242312
rect 317418 241576 317474 241632
rect 345018 241576 345074 241632
rect 350446 242256 350502 242312
rect 373998 241576 374054 241632
rect 378046 242256 378102 242312
rect 405646 242256 405702 242312
rect 401598 241576 401654 241632
rect 434626 242256 434682 242312
rect 429198 241576 429254 241632
rect 462226 242256 462282 242312
rect 458178 241576 458234 241632
rect 489826 242256 489882 242312
rect 485778 241576 485834 241632
rect 238666 215192 238722 215248
rect 238666 188264 238722 188320
rect 266266 215192 266322 215248
rect 262218 214512 262274 214568
rect 293866 215192 293922 215248
rect 289818 214512 289874 214568
rect 322846 215192 322902 215248
rect 317418 214512 317474 214568
rect 345018 214512 345074 214568
rect 350446 215192 350502 215248
rect 373998 214512 374054 214568
rect 378046 215192 378102 215248
rect 405646 215192 405702 215248
rect 401598 214512 401654 214568
rect 434626 215192 434682 215248
rect 429198 214512 429254 214568
rect 462226 215192 462282 215248
rect 458178 214512 458234 214568
rect 489826 215192 489882 215248
rect 485778 214512 485834 214568
rect 266266 188264 266322 188320
rect 262218 187584 262274 187640
rect 293866 188264 293922 188320
rect 289818 187584 289874 187640
rect 322846 188264 322902 188320
rect 317418 187584 317474 187640
rect 345018 187584 345074 187640
rect 350446 188264 350502 188320
rect 373998 187584 374054 187640
rect 378046 188264 378102 188320
rect 405646 188264 405702 188320
rect 401598 187584 401654 187640
rect 434626 188264 434682 188320
rect 429198 187584 429254 187640
rect 462226 188264 462282 188320
rect 458178 187584 458234 187640
rect 489826 188264 489882 188320
rect 485778 187584 485834 187640
rect 238666 161200 238722 161256
rect 266266 161200 266322 161256
rect 262218 160520 262274 160576
rect 293866 161200 293922 161256
rect 289818 160520 289874 160576
rect 322846 161200 322902 161256
rect 317418 160520 317474 160576
rect 345018 160520 345074 160576
rect 350446 161200 350502 161256
rect 373998 160520 374054 160576
rect 378046 161200 378102 161256
rect 405646 161200 405702 161256
rect 401598 160520 401654 160576
rect 434626 161200 434682 161256
rect 429198 160520 429254 160576
rect 462226 161200 462282 161256
rect 458178 160520 458234 160576
rect 489826 161200 489882 161256
rect 485778 160520 485834 160576
rect 238666 134272 238722 134328
rect 266266 134272 266322 134328
rect 262218 133592 262274 133648
rect 293866 134272 293922 134328
rect 289818 133592 289874 133648
rect 322846 134272 322902 134328
rect 317418 133592 317474 133648
rect 345018 133592 345074 133648
rect 350446 134272 350502 134328
rect 373998 133592 374054 133648
rect 378046 134272 378102 134328
rect 405646 134272 405702 134328
rect 401598 133592 401654 133648
rect 434626 134272 434682 134328
rect 429198 133592 429254 133648
rect 462226 134272 462282 134328
rect 458178 133592 458234 133648
rect 489826 134272 489882 134328
rect 485778 133592 485834 133648
rect 238666 107208 238722 107264
rect 238666 80280 238722 80336
rect 266266 107208 266322 107264
rect 262218 106528 262274 106584
rect 293866 107208 293922 107264
rect 289818 106528 289874 106584
rect 322846 107208 322902 107264
rect 317418 106528 317474 106584
rect 345018 106528 345074 106584
rect 350446 107208 350502 107264
rect 373998 106528 374054 106584
rect 378046 107208 378102 107264
rect 405646 107208 405702 107264
rect 401598 106528 401654 106584
rect 434626 107208 434682 107264
rect 429198 106528 429254 106584
rect 462226 107208 462282 107264
rect 458178 106528 458234 106584
rect 489826 107208 489882 107264
rect 485778 106528 485834 106584
rect 266266 80280 266322 80336
rect 262218 79600 262274 79656
rect 293866 80280 293922 80336
rect 289818 79600 289874 79656
rect 322846 80280 322902 80336
rect 317418 79600 317474 79656
rect 345018 79600 345074 79656
rect 350446 80280 350502 80336
rect 373998 79600 374054 79656
rect 378046 80280 378102 80336
rect 405646 80280 405702 80336
rect 401598 79600 401654 79656
rect 434626 80280 434682 80336
rect 429198 79600 429254 79656
rect 462226 80280 462282 80336
rect 458178 79600 458234 79656
rect 489826 80280 489882 80336
rect 485778 79600 485834 79656
rect 238666 53216 238722 53272
rect 70306 26832 70362 26888
rect 97906 26288 97962 26344
rect 93858 25608 93914 25664
rect 121458 25608 121514 25664
rect 126886 26288 126942 26344
rect 154486 26288 154542 26344
rect 149058 25608 149114 25664
rect 178038 25608 178094 25664
rect 182086 26288 182142 26344
rect 209686 26288 209742 26344
rect 205638 25880 205694 25936
rect 238666 26288 238722 26344
rect 233238 25608 233294 25664
rect 266266 53216 266322 53272
rect 262218 52536 262274 52592
rect 293866 53216 293922 53272
rect 289818 52536 289874 52592
rect 322846 53216 322902 53272
rect 317418 52536 317474 52592
rect 345018 52536 345074 52592
rect 350446 53216 350502 53272
rect 373998 52536 374054 52592
rect 378046 53216 378102 53272
rect 405646 53216 405702 53272
rect 401598 52536 401654 52592
rect 434626 53216 434682 53272
rect 429198 52536 429254 52592
rect 462226 53216 462282 53272
rect 458178 52536 458234 52592
rect 489826 53216 489882 53272
rect 485778 52536 485834 52592
rect 266266 26288 266322 26344
rect 262218 25608 262274 25664
rect 293866 26288 293922 26344
rect 289818 25608 289874 25664
rect 317418 25608 317474 25664
rect 322846 26288 322902 26344
rect 345018 25608 345074 25664
rect 350446 26288 350502 26344
rect 373998 25608 374054 25664
rect 378046 26288 378102 26344
rect 405646 26288 405702 26344
rect 401598 25608 401654 25664
rect 434626 26288 434682 26344
rect 429198 25608 429254 25664
rect 462226 26288 462282 26344
rect 458178 25608 458234 25664
rect 489826 26288 489882 26344
rect 485778 25608 485834 25664
rect 518806 674192 518862 674248
rect 513378 673512 513434 673568
rect 518806 647264 518862 647320
rect 513378 646584 513434 646640
rect 518806 620200 518862 620256
rect 513378 619520 513434 619576
rect 518806 593272 518862 593328
rect 513378 592592 513434 592648
rect 518806 566208 518862 566264
rect 513378 565528 513434 565584
rect 518806 539280 518862 539336
rect 513378 538600 513434 538656
rect 518806 512216 518862 512272
rect 513378 511536 513434 511592
rect 540886 510992 540942 511048
rect 518806 485288 518862 485344
rect 513378 484608 513434 484664
rect 518806 458224 518862 458280
rect 513378 457544 513434 457600
rect 518806 431296 518862 431352
rect 513378 430616 513434 430672
rect 518806 404232 518862 404288
rect 513378 403552 513434 403608
rect 518806 377032 518862 377088
rect 513378 375944 513434 376000
rect 540886 375944 540942 376000
rect 518806 350240 518862 350296
rect 513378 349560 513434 349616
rect 518806 322904 518862 322960
rect 513378 322768 513434 322824
rect 518806 296248 518862 296304
rect 513378 295568 513434 295624
rect 518806 269184 518862 269240
rect 513378 268504 513434 268560
rect 518806 242256 518862 242312
rect 513378 241576 513434 241632
rect 518806 215192 518862 215248
rect 513378 214512 513434 214568
rect 518806 188264 518862 188320
rect 513378 187584 513434 187640
rect 518806 161200 518862 161256
rect 513378 160520 513434 160576
rect 518806 134272 518862 134328
rect 513378 133592 513434 133648
rect 518806 107208 518862 107264
rect 513378 106528 513434 106584
rect 518806 80280 518862 80336
rect 513378 79600 513434 79656
rect 518806 53216 518862 53272
rect 513378 52536 513434 52592
rect 513378 25608 513434 25664
rect 518806 26288 518862 26344
rect 542358 673512 542414 673568
rect 545118 674192 545174 674248
rect 569958 673512 570014 673568
rect 542358 646584 542414 646640
rect 545762 647264 545818 647320
rect 542358 619520 542414 619576
rect 545762 620200 545818 620256
rect 542358 592592 542414 592648
rect 545762 593272 545818 593328
rect 542358 565528 542414 565584
rect 545762 566208 545818 566264
rect 542358 538600 542414 538656
rect 545762 539280 545818 539336
rect 545762 512216 545818 512272
rect 542358 484608 542414 484664
rect 545762 485288 545818 485344
rect 542358 457544 542414 457600
rect 545762 458224 545818 458280
rect 542358 430616 542414 430672
rect 545762 431840 545818 431896
rect 542358 403552 542414 403608
rect 545762 404232 545818 404288
rect 545762 377848 545818 377904
rect 542358 349560 542414 349616
rect 545762 350240 545818 350296
rect 542358 321952 542414 322008
rect 545762 323856 545818 323912
rect 542358 295568 542414 295624
rect 545762 296248 545818 296304
rect 542358 268504 542414 268560
rect 545762 269728 545818 269784
rect 542358 241576 542414 241632
rect 545762 242256 545818 242312
rect 542358 214512 542414 214568
rect 545762 215192 545818 215248
rect 542358 187584 542414 187640
rect 545762 188264 545818 188320
rect 542358 160520 542414 160576
rect 545762 161200 545818 161256
rect 542358 133592 542414 133648
rect 545762 134272 545818 134328
rect 542358 106528 542414 106584
rect 545762 107208 545818 107264
rect 542358 79600 542414 79656
rect 545762 80280 545818 80336
rect 542358 52536 542414 52592
rect 545762 53216 545818 53272
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 569958 646584 570014 646640
rect 569958 619520 570014 619576
rect 542358 25608 542414 25664
rect 545762 26288 545818 26344
rect 580170 617480 580226 617536
rect 569958 592592 570014 592648
rect 569958 565528 570014 565584
rect 580262 564304 580318 564360
rect 569958 538600 570014 538656
rect 569958 511536 570014 511592
rect 569958 484608 570014 484664
rect 569958 457544 570014 457600
rect 569958 430616 570014 430672
rect 569958 403552 570014 403608
rect 569958 375944 570014 376000
rect 569958 349560 570014 349616
rect 569958 321952 570014 322008
rect 569958 295568 570014 295624
rect 569958 268504 570014 268560
rect 569958 241576 570014 241632
rect 569958 214512 570014 214568
rect 569958 187584 570014 187640
rect 569958 160520 570014 160576
rect 569958 133592 570014 133648
rect 569958 106528 570014 106584
rect 569958 79600 570014 79656
rect 569958 52536 570014 52592
rect 569958 25608 570014 25664
rect 3422 6432 3478 6488
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 583520 683756 584960 683996
rect 13721 674250 13787 674253
rect 42701 674250 42767 674253
rect 97901 674250 97967 674253
rect 126881 674250 126947 674253
rect 154481 674250 154547 674253
rect 182081 674250 182147 674253
rect 209681 674250 209747 674253
rect 238661 674250 238727 674253
rect 266261 674250 266327 674253
rect 293861 674250 293927 674253
rect 322841 674250 322907 674253
rect 350441 674250 350507 674253
rect 378041 674250 378107 674253
rect 405641 674250 405707 674253
rect 434621 674250 434687 674253
rect 462221 674250 462287 674253
rect 489821 674250 489887 674253
rect 518801 674250 518867 674253
rect 545113 674250 545179 674253
rect 13721 674248 16100 674250
rect 13721 674192 13726 674248
rect 13782 674192 16100 674248
rect 13721 674190 16100 674192
rect 42701 674248 44068 674250
rect 42701 674192 42706 674248
rect 42762 674192 44068 674248
rect 97901 674248 100188 674250
rect 42701 674190 44068 674192
rect 13721 674187 13787 674190
rect 42701 674187 42767 674190
rect 70301 673842 70367 673845
rect 72006 673842 72066 674220
rect 97901 674192 97906 674248
rect 97962 674192 100188 674248
rect 97901 674190 100188 674192
rect 126881 674248 128156 674250
rect 126881 674192 126886 674248
rect 126942 674192 128156 674248
rect 126881 674190 128156 674192
rect 154481 674248 156124 674250
rect 154481 674192 154486 674248
rect 154542 674192 156124 674248
rect 154481 674190 156124 674192
rect 182081 674248 184092 674250
rect 182081 674192 182086 674248
rect 182142 674192 184092 674248
rect 182081 674190 184092 674192
rect 209681 674248 212060 674250
rect 209681 674192 209686 674248
rect 209742 674192 212060 674248
rect 209681 674190 212060 674192
rect 238661 674248 240212 674250
rect 238661 674192 238666 674248
rect 238722 674192 240212 674248
rect 238661 674190 240212 674192
rect 266261 674248 268180 674250
rect 266261 674192 266266 674248
rect 266322 674192 268180 674248
rect 266261 674190 268180 674192
rect 293861 674248 296148 674250
rect 293861 674192 293866 674248
rect 293922 674192 296148 674248
rect 293861 674190 296148 674192
rect 322841 674248 324116 674250
rect 322841 674192 322846 674248
rect 322902 674192 324116 674248
rect 322841 674190 324116 674192
rect 350441 674248 352084 674250
rect 350441 674192 350446 674248
rect 350502 674192 352084 674248
rect 350441 674190 352084 674192
rect 378041 674248 380052 674250
rect 378041 674192 378046 674248
rect 378102 674192 380052 674248
rect 378041 674190 380052 674192
rect 405641 674248 408204 674250
rect 405641 674192 405646 674248
rect 405702 674192 408204 674248
rect 405641 674190 408204 674192
rect 434621 674248 436172 674250
rect 434621 674192 434626 674248
rect 434682 674192 436172 674248
rect 434621 674190 436172 674192
rect 462221 674248 464140 674250
rect 462221 674192 462226 674248
rect 462282 674192 464140 674248
rect 462221 674190 464140 674192
rect 489821 674248 492108 674250
rect 489821 674192 489826 674248
rect 489882 674192 492108 674248
rect 489821 674190 492108 674192
rect 518801 674248 520076 674250
rect 518801 674192 518806 674248
rect 518862 674192 520076 674248
rect 518801 674190 520076 674192
rect 545113 674248 548044 674250
rect 545113 674192 545118 674248
rect 545174 674192 548044 674248
rect 545113 674190 548044 674192
rect 97901 674187 97967 674190
rect 126881 674187 126947 674190
rect 154481 674187 154547 674190
rect 182081 674187 182147 674190
rect 209681 674187 209747 674190
rect 238661 674187 238727 674190
rect 266261 674187 266327 674190
rect 293861 674187 293927 674190
rect 322841 674187 322907 674190
rect 350441 674187 350507 674190
rect 378041 674187 378107 674190
rect 405641 674187 405707 674190
rect 434621 674187 434687 674190
rect 462221 674187 462287 674190
rect 489821 674187 489887 674190
rect 518801 674187 518867 674190
rect 545113 674187 545179 674190
rect 205633 674114 205699 674117
rect 70301 673840 72066 673842
rect 70301 673784 70306 673840
rect 70362 673784 72066 673840
rect 70301 673782 72066 673784
rect 203934 674112 205699 674114
rect 203934 674056 205638 674112
rect 205694 674056 205699 674112
rect 203934 674054 205699 674056
rect 70301 673779 70367 673782
rect 37917 673570 37983 673573
rect 66253 673570 66319 673573
rect 93853 673570 93919 673573
rect 121453 673570 121519 673573
rect 149053 673570 149119 673573
rect 178033 673570 178099 673573
rect 35788 673568 37983 673570
rect 35788 673512 37922 673568
rect 37978 673512 37983 673568
rect 35788 673510 37983 673512
rect 63940 673568 66319 673570
rect 63940 673512 66258 673568
rect 66314 673512 66319 673568
rect 63940 673510 66319 673512
rect 91908 673568 93919 673570
rect 91908 673512 93858 673568
rect 93914 673512 93919 673568
rect 91908 673510 93919 673512
rect 119876 673568 121519 673570
rect 119876 673512 121458 673568
rect 121514 673512 121519 673568
rect 119876 673510 121519 673512
rect 147844 673568 149119 673570
rect 147844 673512 149058 673568
rect 149114 673512 149119 673568
rect 147844 673510 149119 673512
rect 175812 673568 178099 673570
rect 175812 673512 178038 673568
rect 178094 673512 178099 673568
rect 203934 673540 203994 674054
rect 205633 674051 205699 674054
rect 233233 673570 233299 673573
rect 262213 673570 262279 673573
rect 289813 673570 289879 673573
rect 317413 673570 317479 673573
rect 345013 673570 345079 673573
rect 373993 673570 374059 673573
rect 401593 673570 401659 673573
rect 429193 673570 429259 673573
rect 458173 673570 458239 673573
rect 485773 673570 485839 673573
rect 513373 673570 513439 673573
rect 542353 673570 542419 673573
rect 569953 673570 570019 673573
rect 231932 673568 233299 673570
rect 175812 673510 178099 673512
rect 231932 673512 233238 673568
rect 233294 673512 233299 673568
rect 231932 673510 233299 673512
rect 259900 673568 262279 673570
rect 259900 673512 262218 673568
rect 262274 673512 262279 673568
rect 259900 673510 262279 673512
rect 287868 673568 289879 673570
rect 287868 673512 289818 673568
rect 289874 673512 289879 673568
rect 287868 673510 289879 673512
rect 315836 673568 317479 673570
rect 315836 673512 317418 673568
rect 317474 673512 317479 673568
rect 315836 673510 317479 673512
rect 343804 673568 345079 673570
rect 343804 673512 345018 673568
rect 345074 673512 345079 673568
rect 343804 673510 345079 673512
rect 371956 673568 374059 673570
rect 371956 673512 373998 673568
rect 374054 673512 374059 673568
rect 371956 673510 374059 673512
rect 399924 673568 401659 673570
rect 399924 673512 401598 673568
rect 401654 673512 401659 673568
rect 399924 673510 401659 673512
rect 427892 673568 429259 673570
rect 427892 673512 429198 673568
rect 429254 673512 429259 673568
rect 427892 673510 429259 673512
rect 455860 673568 458239 673570
rect 455860 673512 458178 673568
rect 458234 673512 458239 673568
rect 455860 673510 458239 673512
rect 483828 673568 485839 673570
rect 483828 673512 485778 673568
rect 485834 673512 485839 673568
rect 483828 673510 485839 673512
rect 511796 673568 513439 673570
rect 511796 673512 513378 673568
rect 513434 673512 513439 673568
rect 511796 673510 513439 673512
rect 539948 673568 542419 673570
rect 539948 673512 542358 673568
rect 542414 673512 542419 673568
rect 539948 673510 542419 673512
rect 567916 673568 570019 673570
rect 567916 673512 569958 673568
rect 570014 673512 570019 673568
rect 567916 673510 570019 673512
rect 37917 673507 37983 673510
rect 66253 673507 66319 673510
rect 93853 673507 93919 673510
rect 121453 673507 121519 673510
rect 149053 673507 149119 673510
rect 178033 673507 178099 673510
rect 233233 673507 233299 673510
rect 262213 673507 262279 673510
rect 289813 673507 289879 673510
rect 317413 673507 317479 673510
rect 345013 673507 345079 673510
rect 373993 673507 374059 673510
rect 401593 673507 401659 673510
rect 429193 673507 429259 673510
rect 458173 673507 458239 673510
rect 485773 673507 485839 673510
rect 513373 673507 513439 673510
rect 542353 673507 542419 673510
rect 569953 673507 570019 673510
rect -960 671108 480 671348
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect 13721 647322 13787 647325
rect 42701 647322 42767 647325
rect 70301 647322 70367 647325
rect 97901 647322 97967 647325
rect 126881 647322 126947 647325
rect 154481 647322 154547 647325
rect 182081 647322 182147 647325
rect 209681 647322 209747 647325
rect 238661 647322 238727 647325
rect 266261 647322 266327 647325
rect 293861 647322 293927 647325
rect 322841 647322 322907 647325
rect 350441 647322 350507 647325
rect 378041 647322 378107 647325
rect 405641 647322 405707 647325
rect 434621 647322 434687 647325
rect 462221 647322 462287 647325
rect 489821 647322 489887 647325
rect 518801 647322 518867 647325
rect 545757 647322 545823 647325
rect 13721 647320 16100 647322
rect 13721 647264 13726 647320
rect 13782 647264 16100 647320
rect 13721 647262 16100 647264
rect 42701 647320 44068 647322
rect 42701 647264 42706 647320
rect 42762 647264 44068 647320
rect 42701 647262 44068 647264
rect 70301 647320 72036 647322
rect 70301 647264 70306 647320
rect 70362 647264 72036 647320
rect 70301 647262 72036 647264
rect 97901 647320 100188 647322
rect 97901 647264 97906 647320
rect 97962 647264 100188 647320
rect 97901 647262 100188 647264
rect 126881 647320 128156 647322
rect 126881 647264 126886 647320
rect 126942 647264 128156 647320
rect 126881 647262 128156 647264
rect 154481 647320 156124 647322
rect 154481 647264 154486 647320
rect 154542 647264 156124 647320
rect 154481 647262 156124 647264
rect 182081 647320 184092 647322
rect 182081 647264 182086 647320
rect 182142 647264 184092 647320
rect 182081 647262 184092 647264
rect 209681 647320 212060 647322
rect 209681 647264 209686 647320
rect 209742 647264 212060 647320
rect 209681 647262 212060 647264
rect 238661 647320 240212 647322
rect 238661 647264 238666 647320
rect 238722 647264 240212 647320
rect 238661 647262 240212 647264
rect 266261 647320 268180 647322
rect 266261 647264 266266 647320
rect 266322 647264 268180 647320
rect 266261 647262 268180 647264
rect 293861 647320 296148 647322
rect 293861 647264 293866 647320
rect 293922 647264 296148 647320
rect 293861 647262 296148 647264
rect 322841 647320 324116 647322
rect 322841 647264 322846 647320
rect 322902 647264 324116 647320
rect 322841 647262 324116 647264
rect 350441 647320 352084 647322
rect 350441 647264 350446 647320
rect 350502 647264 352084 647320
rect 350441 647262 352084 647264
rect 378041 647320 380052 647322
rect 378041 647264 378046 647320
rect 378102 647264 380052 647320
rect 378041 647262 380052 647264
rect 405641 647320 408204 647322
rect 405641 647264 405646 647320
rect 405702 647264 408204 647320
rect 405641 647262 408204 647264
rect 434621 647320 436172 647322
rect 434621 647264 434626 647320
rect 434682 647264 436172 647320
rect 434621 647262 436172 647264
rect 462221 647320 464140 647322
rect 462221 647264 462226 647320
rect 462282 647264 464140 647320
rect 462221 647262 464140 647264
rect 489821 647320 492108 647322
rect 489821 647264 489826 647320
rect 489882 647264 492108 647320
rect 489821 647262 492108 647264
rect 518801 647320 520076 647322
rect 518801 647264 518806 647320
rect 518862 647264 520076 647320
rect 518801 647262 520076 647264
rect 545757 647320 548044 647322
rect 545757 647264 545762 647320
rect 545818 647264 548044 647320
rect 545757 647262 548044 647264
rect 13721 647259 13787 647262
rect 42701 647259 42767 647262
rect 70301 647259 70367 647262
rect 97901 647259 97967 647262
rect 126881 647259 126947 647262
rect 154481 647259 154547 647262
rect 182081 647259 182147 647262
rect 209681 647259 209747 647262
rect 238661 647259 238727 647262
rect 266261 647259 266327 647262
rect 293861 647259 293927 647262
rect 322841 647259 322907 647262
rect 350441 647259 350507 647262
rect 378041 647259 378107 647262
rect 405641 647259 405707 647262
rect 434621 647259 434687 647262
rect 462221 647259 462287 647262
rect 489821 647259 489887 647262
rect 518801 647259 518867 647262
rect 545757 647259 545823 647262
rect 37917 646642 37983 646645
rect 66253 646642 66319 646645
rect 93853 646642 93919 646645
rect 121453 646642 121519 646645
rect 149053 646642 149119 646645
rect 178033 646642 178099 646645
rect 205633 646642 205699 646645
rect 233233 646642 233299 646645
rect 262213 646642 262279 646645
rect 289813 646642 289879 646645
rect 317413 646642 317479 646645
rect 345013 646642 345079 646645
rect 373993 646642 374059 646645
rect 401593 646642 401659 646645
rect 429193 646642 429259 646645
rect 458173 646642 458239 646645
rect 485773 646642 485839 646645
rect 513373 646642 513439 646645
rect 542353 646642 542419 646645
rect 569953 646642 570019 646645
rect 35788 646640 37983 646642
rect 35788 646584 37922 646640
rect 37978 646584 37983 646640
rect 35788 646582 37983 646584
rect 63940 646640 66319 646642
rect 63940 646584 66258 646640
rect 66314 646584 66319 646640
rect 63940 646582 66319 646584
rect 91908 646640 93919 646642
rect 91908 646584 93858 646640
rect 93914 646584 93919 646640
rect 91908 646582 93919 646584
rect 119876 646640 121519 646642
rect 119876 646584 121458 646640
rect 121514 646584 121519 646640
rect 119876 646582 121519 646584
rect 147844 646640 149119 646642
rect 147844 646584 149058 646640
rect 149114 646584 149119 646640
rect 147844 646582 149119 646584
rect 175812 646640 178099 646642
rect 175812 646584 178038 646640
rect 178094 646584 178099 646640
rect 175812 646582 178099 646584
rect 203964 646640 205699 646642
rect 203964 646584 205638 646640
rect 205694 646584 205699 646640
rect 203964 646582 205699 646584
rect 231932 646640 233299 646642
rect 231932 646584 233238 646640
rect 233294 646584 233299 646640
rect 231932 646582 233299 646584
rect 259900 646640 262279 646642
rect 259900 646584 262218 646640
rect 262274 646584 262279 646640
rect 259900 646582 262279 646584
rect 287868 646640 289879 646642
rect 287868 646584 289818 646640
rect 289874 646584 289879 646640
rect 287868 646582 289879 646584
rect 315836 646640 317479 646642
rect 315836 646584 317418 646640
rect 317474 646584 317479 646640
rect 315836 646582 317479 646584
rect 343804 646640 345079 646642
rect 343804 646584 345018 646640
rect 345074 646584 345079 646640
rect 343804 646582 345079 646584
rect 371956 646640 374059 646642
rect 371956 646584 373998 646640
rect 374054 646584 374059 646640
rect 371956 646582 374059 646584
rect 399924 646640 401659 646642
rect 399924 646584 401598 646640
rect 401654 646584 401659 646640
rect 399924 646582 401659 646584
rect 427892 646640 429259 646642
rect 427892 646584 429198 646640
rect 429254 646584 429259 646640
rect 427892 646582 429259 646584
rect 455860 646640 458239 646642
rect 455860 646584 458178 646640
rect 458234 646584 458239 646640
rect 455860 646582 458239 646584
rect 483828 646640 485839 646642
rect 483828 646584 485778 646640
rect 485834 646584 485839 646640
rect 483828 646582 485839 646584
rect 511796 646640 513439 646642
rect 511796 646584 513378 646640
rect 513434 646584 513439 646640
rect 511796 646582 513439 646584
rect 539948 646640 542419 646642
rect 539948 646584 542358 646640
rect 542414 646584 542419 646640
rect 539948 646582 542419 646584
rect 567916 646640 570019 646642
rect 567916 646584 569958 646640
rect 570014 646584 570019 646640
rect 567916 646582 570019 646584
rect 37917 646579 37983 646582
rect 66253 646579 66319 646582
rect 93853 646579 93919 646582
rect 121453 646579 121519 646582
rect 149053 646579 149119 646582
rect 178033 646579 178099 646582
rect 205633 646579 205699 646582
rect 233233 646579 233299 646582
rect 262213 646579 262279 646582
rect 289813 646579 289879 646582
rect 317413 646579 317479 646582
rect 345013 646579 345079 646582
rect 373993 646579 374059 646582
rect 401593 646579 401659 646582
rect 429193 646579 429259 646582
rect 458173 646579 458239 646582
rect 485773 646579 485839 646582
rect 513373 646579 513439 646582
rect 542353 646579 542419 646582
rect 569953 646579 570019 646582
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 632090 480 632180
rect 3141 632090 3207 632093
rect -960 632088 3207 632090
rect -960 632032 3146 632088
rect 3202 632032 3207 632088
rect -960 632030 3207 632032
rect -960 631940 480 632030
rect 3141 632027 3207 632030
rect 583520 630716 584960 630956
rect 13721 620258 13787 620261
rect 42701 620258 42767 620261
rect 70301 620258 70367 620261
rect 97901 620258 97967 620261
rect 126881 620258 126947 620261
rect 154481 620258 154547 620261
rect 182081 620258 182147 620261
rect 209681 620258 209747 620261
rect 238661 620258 238727 620261
rect 266261 620258 266327 620261
rect 293861 620258 293927 620261
rect 322841 620258 322907 620261
rect 350441 620258 350507 620261
rect 378041 620258 378107 620261
rect 405641 620258 405707 620261
rect 434621 620258 434687 620261
rect 462221 620258 462287 620261
rect 489821 620258 489887 620261
rect 518801 620258 518867 620261
rect 545757 620258 545823 620261
rect 13721 620256 16100 620258
rect 13721 620200 13726 620256
rect 13782 620200 16100 620256
rect 13721 620198 16100 620200
rect 42701 620256 44068 620258
rect 42701 620200 42706 620256
rect 42762 620200 44068 620256
rect 42701 620198 44068 620200
rect 70301 620256 72036 620258
rect 70301 620200 70306 620256
rect 70362 620200 72036 620256
rect 70301 620198 72036 620200
rect 97901 620256 100188 620258
rect 97901 620200 97906 620256
rect 97962 620200 100188 620256
rect 97901 620198 100188 620200
rect 126881 620256 128156 620258
rect 126881 620200 126886 620256
rect 126942 620200 128156 620256
rect 126881 620198 128156 620200
rect 154481 620256 156124 620258
rect 154481 620200 154486 620256
rect 154542 620200 156124 620256
rect 154481 620198 156124 620200
rect 182081 620256 184092 620258
rect 182081 620200 182086 620256
rect 182142 620200 184092 620256
rect 182081 620198 184092 620200
rect 209681 620256 212060 620258
rect 209681 620200 209686 620256
rect 209742 620200 212060 620256
rect 209681 620198 212060 620200
rect 238661 620256 240212 620258
rect 238661 620200 238666 620256
rect 238722 620200 240212 620256
rect 238661 620198 240212 620200
rect 266261 620256 268180 620258
rect 266261 620200 266266 620256
rect 266322 620200 268180 620256
rect 266261 620198 268180 620200
rect 293861 620256 296148 620258
rect 293861 620200 293866 620256
rect 293922 620200 296148 620256
rect 293861 620198 296148 620200
rect 322841 620256 324116 620258
rect 322841 620200 322846 620256
rect 322902 620200 324116 620256
rect 322841 620198 324116 620200
rect 350441 620256 352084 620258
rect 350441 620200 350446 620256
rect 350502 620200 352084 620256
rect 350441 620198 352084 620200
rect 378041 620256 380052 620258
rect 378041 620200 378046 620256
rect 378102 620200 380052 620256
rect 378041 620198 380052 620200
rect 405641 620256 408204 620258
rect 405641 620200 405646 620256
rect 405702 620200 408204 620256
rect 405641 620198 408204 620200
rect 434621 620256 436172 620258
rect 434621 620200 434626 620256
rect 434682 620200 436172 620256
rect 434621 620198 436172 620200
rect 462221 620256 464140 620258
rect 462221 620200 462226 620256
rect 462282 620200 464140 620256
rect 462221 620198 464140 620200
rect 489821 620256 492108 620258
rect 489821 620200 489826 620256
rect 489882 620200 492108 620256
rect 489821 620198 492108 620200
rect 518801 620256 520076 620258
rect 518801 620200 518806 620256
rect 518862 620200 520076 620256
rect 518801 620198 520076 620200
rect 545757 620256 548044 620258
rect 545757 620200 545762 620256
rect 545818 620200 548044 620256
rect 545757 620198 548044 620200
rect 13721 620195 13787 620198
rect 42701 620195 42767 620198
rect 70301 620195 70367 620198
rect 97901 620195 97967 620198
rect 126881 620195 126947 620198
rect 154481 620195 154547 620198
rect 182081 620195 182147 620198
rect 209681 620195 209747 620198
rect 238661 620195 238727 620198
rect 266261 620195 266327 620198
rect 293861 620195 293927 620198
rect 322841 620195 322907 620198
rect 350441 620195 350507 620198
rect 378041 620195 378107 620198
rect 405641 620195 405707 620198
rect 434621 620195 434687 620198
rect 462221 620195 462287 620198
rect 489821 620195 489887 620198
rect 518801 620195 518867 620198
rect 545757 620195 545823 620198
rect 37917 619578 37983 619581
rect 66253 619578 66319 619581
rect 93853 619578 93919 619581
rect 121453 619578 121519 619581
rect 149053 619578 149119 619581
rect 178033 619578 178099 619581
rect 205633 619578 205699 619581
rect 233233 619578 233299 619581
rect 262213 619578 262279 619581
rect 289813 619578 289879 619581
rect 317413 619578 317479 619581
rect 345013 619578 345079 619581
rect 373993 619578 374059 619581
rect 401593 619578 401659 619581
rect 429193 619578 429259 619581
rect 458173 619578 458239 619581
rect 485773 619578 485839 619581
rect 513373 619578 513439 619581
rect 542353 619578 542419 619581
rect 569953 619578 570019 619581
rect 35788 619576 37983 619578
rect 35788 619520 37922 619576
rect 37978 619520 37983 619576
rect 35788 619518 37983 619520
rect 63940 619576 66319 619578
rect 63940 619520 66258 619576
rect 66314 619520 66319 619576
rect 63940 619518 66319 619520
rect 91908 619576 93919 619578
rect 91908 619520 93858 619576
rect 93914 619520 93919 619576
rect 91908 619518 93919 619520
rect 119876 619576 121519 619578
rect 119876 619520 121458 619576
rect 121514 619520 121519 619576
rect 119876 619518 121519 619520
rect 147844 619576 149119 619578
rect 147844 619520 149058 619576
rect 149114 619520 149119 619576
rect 147844 619518 149119 619520
rect 175812 619576 178099 619578
rect 175812 619520 178038 619576
rect 178094 619520 178099 619576
rect 175812 619518 178099 619520
rect 203964 619576 205699 619578
rect 203964 619520 205638 619576
rect 205694 619520 205699 619576
rect 203964 619518 205699 619520
rect 231932 619576 233299 619578
rect 231932 619520 233238 619576
rect 233294 619520 233299 619576
rect 231932 619518 233299 619520
rect 259900 619576 262279 619578
rect 259900 619520 262218 619576
rect 262274 619520 262279 619576
rect 259900 619518 262279 619520
rect 287868 619576 289879 619578
rect 287868 619520 289818 619576
rect 289874 619520 289879 619576
rect 287868 619518 289879 619520
rect 315836 619576 317479 619578
rect 315836 619520 317418 619576
rect 317474 619520 317479 619576
rect 315836 619518 317479 619520
rect 343804 619576 345079 619578
rect 343804 619520 345018 619576
rect 345074 619520 345079 619576
rect 343804 619518 345079 619520
rect 371956 619576 374059 619578
rect 371956 619520 373998 619576
rect 374054 619520 374059 619576
rect 371956 619518 374059 619520
rect 399924 619576 401659 619578
rect 399924 619520 401598 619576
rect 401654 619520 401659 619576
rect 399924 619518 401659 619520
rect 427892 619576 429259 619578
rect 427892 619520 429198 619576
rect 429254 619520 429259 619576
rect 427892 619518 429259 619520
rect 455860 619576 458239 619578
rect 455860 619520 458178 619576
rect 458234 619520 458239 619576
rect 455860 619518 458239 619520
rect 483828 619576 485839 619578
rect 483828 619520 485778 619576
rect 485834 619520 485839 619576
rect 483828 619518 485839 619520
rect 511796 619576 513439 619578
rect 511796 619520 513378 619576
rect 513434 619520 513439 619576
rect 511796 619518 513439 619520
rect 539948 619576 542419 619578
rect 539948 619520 542358 619576
rect 542414 619520 542419 619576
rect 539948 619518 542419 619520
rect 567916 619576 570019 619578
rect 567916 619520 569958 619576
rect 570014 619520 570019 619576
rect 567916 619518 570019 619520
rect 37917 619515 37983 619518
rect 66253 619515 66319 619518
rect 93853 619515 93919 619518
rect 121453 619515 121519 619518
rect 149053 619515 149119 619518
rect 178033 619515 178099 619518
rect 205633 619515 205699 619518
rect 233233 619515 233299 619518
rect 262213 619515 262279 619518
rect 289813 619515 289879 619518
rect 317413 619515 317479 619518
rect 345013 619515 345079 619518
rect 373993 619515 374059 619518
rect 401593 619515 401659 619518
rect 429193 619515 429259 619518
rect 458173 619515 458239 619518
rect 485773 619515 485839 619518
rect 513373 619515 513439 619518
rect 542353 619515 542419 619518
rect 569953 619515 570019 619518
rect -960 619020 480 619260
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect 13721 593330 13787 593333
rect 42701 593330 42767 593333
rect 70301 593330 70367 593333
rect 97901 593330 97967 593333
rect 126881 593330 126947 593333
rect 154481 593330 154547 593333
rect 182081 593330 182147 593333
rect 209681 593330 209747 593333
rect 238661 593330 238727 593333
rect 266261 593330 266327 593333
rect 293861 593330 293927 593333
rect 322841 593330 322907 593333
rect 350441 593330 350507 593333
rect 378041 593330 378107 593333
rect 405641 593330 405707 593333
rect 434621 593330 434687 593333
rect 462221 593330 462287 593333
rect 489821 593330 489887 593333
rect 518801 593330 518867 593333
rect 545757 593330 545823 593333
rect 13721 593328 16100 593330
rect 13721 593272 13726 593328
rect 13782 593272 16100 593328
rect 13721 593270 16100 593272
rect 42701 593328 44068 593330
rect 42701 593272 42706 593328
rect 42762 593272 44068 593328
rect 42701 593270 44068 593272
rect 70301 593328 72036 593330
rect 70301 593272 70306 593328
rect 70362 593272 72036 593328
rect 70301 593270 72036 593272
rect 97901 593328 100188 593330
rect 97901 593272 97906 593328
rect 97962 593272 100188 593328
rect 97901 593270 100188 593272
rect 126881 593328 128156 593330
rect 126881 593272 126886 593328
rect 126942 593272 128156 593328
rect 126881 593270 128156 593272
rect 154481 593328 156124 593330
rect 154481 593272 154486 593328
rect 154542 593272 156124 593328
rect 154481 593270 156124 593272
rect 182081 593328 184092 593330
rect 182081 593272 182086 593328
rect 182142 593272 184092 593328
rect 182081 593270 184092 593272
rect 209681 593328 212060 593330
rect 209681 593272 209686 593328
rect 209742 593272 212060 593328
rect 209681 593270 212060 593272
rect 238661 593328 240212 593330
rect 238661 593272 238666 593328
rect 238722 593272 240212 593328
rect 238661 593270 240212 593272
rect 266261 593328 268180 593330
rect 266261 593272 266266 593328
rect 266322 593272 268180 593328
rect 266261 593270 268180 593272
rect 293861 593328 296148 593330
rect 293861 593272 293866 593328
rect 293922 593272 296148 593328
rect 293861 593270 296148 593272
rect 322841 593328 324116 593330
rect 322841 593272 322846 593328
rect 322902 593272 324116 593328
rect 322841 593270 324116 593272
rect 350441 593328 352084 593330
rect 350441 593272 350446 593328
rect 350502 593272 352084 593328
rect 350441 593270 352084 593272
rect 378041 593328 380052 593330
rect 378041 593272 378046 593328
rect 378102 593272 380052 593328
rect 378041 593270 380052 593272
rect 405641 593328 408204 593330
rect 405641 593272 405646 593328
rect 405702 593272 408204 593328
rect 405641 593270 408204 593272
rect 434621 593328 436172 593330
rect 434621 593272 434626 593328
rect 434682 593272 436172 593328
rect 434621 593270 436172 593272
rect 462221 593328 464140 593330
rect 462221 593272 462226 593328
rect 462282 593272 464140 593328
rect 462221 593270 464140 593272
rect 489821 593328 492108 593330
rect 489821 593272 489826 593328
rect 489882 593272 492108 593328
rect 489821 593270 492108 593272
rect 518801 593328 520076 593330
rect 518801 593272 518806 593328
rect 518862 593272 520076 593328
rect 518801 593270 520076 593272
rect 545757 593328 548044 593330
rect 545757 593272 545762 593328
rect 545818 593272 548044 593328
rect 545757 593270 548044 593272
rect 13721 593267 13787 593270
rect 42701 593267 42767 593270
rect 70301 593267 70367 593270
rect 97901 593267 97967 593270
rect 126881 593267 126947 593270
rect 154481 593267 154547 593270
rect 182081 593267 182147 593270
rect 209681 593267 209747 593270
rect 238661 593267 238727 593270
rect 266261 593267 266327 593270
rect 293861 593267 293927 593270
rect 322841 593267 322907 593270
rect 350441 593267 350507 593270
rect 378041 593267 378107 593270
rect 405641 593267 405707 593270
rect 434621 593267 434687 593270
rect 462221 593267 462287 593270
rect 489821 593267 489887 593270
rect 518801 593267 518867 593270
rect 545757 593267 545823 593270
rect -960 592908 480 593148
rect 37917 592650 37983 592653
rect 66253 592650 66319 592653
rect 93853 592650 93919 592653
rect 121453 592650 121519 592653
rect 149053 592650 149119 592653
rect 178033 592650 178099 592653
rect 205633 592650 205699 592653
rect 233233 592650 233299 592653
rect 262213 592650 262279 592653
rect 289813 592650 289879 592653
rect 317413 592650 317479 592653
rect 345013 592650 345079 592653
rect 373993 592650 374059 592653
rect 401593 592650 401659 592653
rect 429193 592650 429259 592653
rect 458173 592650 458239 592653
rect 485773 592650 485839 592653
rect 513373 592650 513439 592653
rect 542353 592650 542419 592653
rect 569953 592650 570019 592653
rect 35788 592648 37983 592650
rect 35788 592592 37922 592648
rect 37978 592592 37983 592648
rect 35788 592590 37983 592592
rect 63940 592648 66319 592650
rect 63940 592592 66258 592648
rect 66314 592592 66319 592648
rect 63940 592590 66319 592592
rect 91908 592648 93919 592650
rect 91908 592592 93858 592648
rect 93914 592592 93919 592648
rect 91908 592590 93919 592592
rect 119876 592648 121519 592650
rect 119876 592592 121458 592648
rect 121514 592592 121519 592648
rect 119876 592590 121519 592592
rect 147844 592648 149119 592650
rect 147844 592592 149058 592648
rect 149114 592592 149119 592648
rect 147844 592590 149119 592592
rect 175812 592648 178099 592650
rect 175812 592592 178038 592648
rect 178094 592592 178099 592648
rect 175812 592590 178099 592592
rect 203964 592648 205699 592650
rect 203964 592592 205638 592648
rect 205694 592592 205699 592648
rect 203964 592590 205699 592592
rect 231932 592648 233299 592650
rect 231932 592592 233238 592648
rect 233294 592592 233299 592648
rect 231932 592590 233299 592592
rect 259900 592648 262279 592650
rect 259900 592592 262218 592648
rect 262274 592592 262279 592648
rect 259900 592590 262279 592592
rect 287868 592648 289879 592650
rect 287868 592592 289818 592648
rect 289874 592592 289879 592648
rect 287868 592590 289879 592592
rect 315836 592648 317479 592650
rect 315836 592592 317418 592648
rect 317474 592592 317479 592648
rect 315836 592590 317479 592592
rect 343804 592648 345079 592650
rect 343804 592592 345018 592648
rect 345074 592592 345079 592648
rect 343804 592590 345079 592592
rect 371956 592648 374059 592650
rect 371956 592592 373998 592648
rect 374054 592592 374059 592648
rect 371956 592590 374059 592592
rect 399924 592648 401659 592650
rect 399924 592592 401598 592648
rect 401654 592592 401659 592648
rect 399924 592590 401659 592592
rect 427892 592648 429259 592650
rect 427892 592592 429198 592648
rect 429254 592592 429259 592648
rect 427892 592590 429259 592592
rect 455860 592648 458239 592650
rect 455860 592592 458178 592648
rect 458234 592592 458239 592648
rect 455860 592590 458239 592592
rect 483828 592648 485839 592650
rect 483828 592592 485778 592648
rect 485834 592592 485839 592648
rect 483828 592590 485839 592592
rect 511796 592648 513439 592650
rect 511796 592592 513378 592648
rect 513434 592592 513439 592648
rect 511796 592590 513439 592592
rect 539948 592648 542419 592650
rect 539948 592592 542358 592648
rect 542414 592592 542419 592648
rect 539948 592590 542419 592592
rect 567916 592648 570019 592650
rect 567916 592592 569958 592648
rect 570014 592592 570019 592648
rect 567916 592590 570019 592592
rect 37917 592587 37983 592590
rect 66253 592587 66319 592590
rect 93853 592587 93919 592590
rect 121453 592587 121519 592590
rect 149053 592587 149119 592590
rect 178033 592587 178099 592590
rect 205633 592587 205699 592590
rect 233233 592587 233299 592590
rect 262213 592587 262279 592590
rect 289813 592587 289879 592590
rect 317413 592587 317479 592590
rect 345013 592587 345079 592590
rect 373993 592587 374059 592590
rect 401593 592587 401659 592590
rect 429193 592587 429259 592590
rect 458173 592587 458239 592590
rect 485773 592587 485839 592590
rect 513373 592587 513439 592590
rect 542353 592587 542419 592590
rect 569953 592587 570019 592590
rect 583520 590868 584960 591108
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 13721 566266 13787 566269
rect 42701 566266 42767 566269
rect 70301 566266 70367 566269
rect 97901 566266 97967 566269
rect 126881 566266 126947 566269
rect 154481 566266 154547 566269
rect 182081 566266 182147 566269
rect 209681 566266 209747 566269
rect 238661 566266 238727 566269
rect 266261 566266 266327 566269
rect 293861 566266 293927 566269
rect 322841 566266 322907 566269
rect 350441 566266 350507 566269
rect 378041 566266 378107 566269
rect 405641 566266 405707 566269
rect 434621 566266 434687 566269
rect 462221 566266 462287 566269
rect 489821 566266 489887 566269
rect 518801 566266 518867 566269
rect 545757 566266 545823 566269
rect 13721 566264 16100 566266
rect 13721 566208 13726 566264
rect 13782 566208 16100 566264
rect 13721 566206 16100 566208
rect 42701 566264 44068 566266
rect 42701 566208 42706 566264
rect 42762 566208 44068 566264
rect 42701 566206 44068 566208
rect 70301 566264 72036 566266
rect 70301 566208 70306 566264
rect 70362 566208 72036 566264
rect 70301 566206 72036 566208
rect 97901 566264 100188 566266
rect 97901 566208 97906 566264
rect 97962 566208 100188 566264
rect 97901 566206 100188 566208
rect 126881 566264 128156 566266
rect 126881 566208 126886 566264
rect 126942 566208 128156 566264
rect 126881 566206 128156 566208
rect 154481 566264 156124 566266
rect 154481 566208 154486 566264
rect 154542 566208 156124 566264
rect 154481 566206 156124 566208
rect 182081 566264 184092 566266
rect 182081 566208 182086 566264
rect 182142 566208 184092 566264
rect 182081 566206 184092 566208
rect 209681 566264 212060 566266
rect 209681 566208 209686 566264
rect 209742 566208 212060 566264
rect 209681 566206 212060 566208
rect 238661 566264 240212 566266
rect 238661 566208 238666 566264
rect 238722 566208 240212 566264
rect 238661 566206 240212 566208
rect 266261 566264 268180 566266
rect 266261 566208 266266 566264
rect 266322 566208 268180 566264
rect 266261 566206 268180 566208
rect 293861 566264 296148 566266
rect 293861 566208 293866 566264
rect 293922 566208 296148 566264
rect 293861 566206 296148 566208
rect 322841 566264 324116 566266
rect 322841 566208 322846 566264
rect 322902 566208 324116 566264
rect 322841 566206 324116 566208
rect 350441 566264 352084 566266
rect 350441 566208 350446 566264
rect 350502 566208 352084 566264
rect 350441 566206 352084 566208
rect 378041 566264 380052 566266
rect 378041 566208 378046 566264
rect 378102 566208 380052 566264
rect 378041 566206 380052 566208
rect 405641 566264 408204 566266
rect 405641 566208 405646 566264
rect 405702 566208 408204 566264
rect 405641 566206 408204 566208
rect 434621 566264 436172 566266
rect 434621 566208 434626 566264
rect 434682 566208 436172 566264
rect 434621 566206 436172 566208
rect 462221 566264 464140 566266
rect 462221 566208 462226 566264
rect 462282 566208 464140 566264
rect 462221 566206 464140 566208
rect 489821 566264 492108 566266
rect 489821 566208 489826 566264
rect 489882 566208 492108 566264
rect 489821 566206 492108 566208
rect 518801 566264 520076 566266
rect 518801 566208 518806 566264
rect 518862 566208 520076 566264
rect 518801 566206 520076 566208
rect 545757 566264 548044 566266
rect 545757 566208 545762 566264
rect 545818 566208 548044 566264
rect 545757 566206 548044 566208
rect 13721 566203 13787 566206
rect 42701 566203 42767 566206
rect 70301 566203 70367 566206
rect 97901 566203 97967 566206
rect 126881 566203 126947 566206
rect 154481 566203 154547 566206
rect 182081 566203 182147 566206
rect 209681 566203 209747 566206
rect 238661 566203 238727 566206
rect 266261 566203 266327 566206
rect 293861 566203 293927 566206
rect 322841 566203 322907 566206
rect 350441 566203 350507 566206
rect 378041 566203 378107 566206
rect 405641 566203 405707 566206
rect 434621 566203 434687 566206
rect 462221 566203 462287 566206
rect 489821 566203 489887 566206
rect 518801 566203 518867 566206
rect 545757 566203 545823 566206
rect 37917 565586 37983 565589
rect 66253 565586 66319 565589
rect 93853 565586 93919 565589
rect 121453 565586 121519 565589
rect 149053 565586 149119 565589
rect 178033 565586 178099 565589
rect 205633 565586 205699 565589
rect 233233 565586 233299 565589
rect 262213 565586 262279 565589
rect 289813 565586 289879 565589
rect 317413 565586 317479 565589
rect 345013 565586 345079 565589
rect 373993 565586 374059 565589
rect 401593 565586 401659 565589
rect 429193 565586 429259 565589
rect 458173 565586 458239 565589
rect 485773 565586 485839 565589
rect 513373 565586 513439 565589
rect 542353 565586 542419 565589
rect 569953 565586 570019 565589
rect 35788 565584 37983 565586
rect 35788 565528 37922 565584
rect 37978 565528 37983 565584
rect 35788 565526 37983 565528
rect 63940 565584 66319 565586
rect 63940 565528 66258 565584
rect 66314 565528 66319 565584
rect 63940 565526 66319 565528
rect 91908 565584 93919 565586
rect 91908 565528 93858 565584
rect 93914 565528 93919 565584
rect 91908 565526 93919 565528
rect 119876 565584 121519 565586
rect 119876 565528 121458 565584
rect 121514 565528 121519 565584
rect 119876 565526 121519 565528
rect 147844 565584 149119 565586
rect 147844 565528 149058 565584
rect 149114 565528 149119 565584
rect 147844 565526 149119 565528
rect 175812 565584 178099 565586
rect 175812 565528 178038 565584
rect 178094 565528 178099 565584
rect 175812 565526 178099 565528
rect 203964 565584 205699 565586
rect 203964 565528 205638 565584
rect 205694 565528 205699 565584
rect 203964 565526 205699 565528
rect 231932 565584 233299 565586
rect 231932 565528 233238 565584
rect 233294 565528 233299 565584
rect 231932 565526 233299 565528
rect 259900 565584 262279 565586
rect 259900 565528 262218 565584
rect 262274 565528 262279 565584
rect 259900 565526 262279 565528
rect 287868 565584 289879 565586
rect 287868 565528 289818 565584
rect 289874 565528 289879 565584
rect 287868 565526 289879 565528
rect 315836 565584 317479 565586
rect 315836 565528 317418 565584
rect 317474 565528 317479 565584
rect 315836 565526 317479 565528
rect 343804 565584 345079 565586
rect 343804 565528 345018 565584
rect 345074 565528 345079 565584
rect 343804 565526 345079 565528
rect 371956 565584 374059 565586
rect 371956 565528 373998 565584
rect 374054 565528 374059 565584
rect 371956 565526 374059 565528
rect 399924 565584 401659 565586
rect 399924 565528 401598 565584
rect 401654 565528 401659 565584
rect 399924 565526 401659 565528
rect 427892 565584 429259 565586
rect 427892 565528 429198 565584
rect 429254 565528 429259 565584
rect 427892 565526 429259 565528
rect 455860 565584 458239 565586
rect 455860 565528 458178 565584
rect 458234 565528 458239 565584
rect 455860 565526 458239 565528
rect 483828 565584 485839 565586
rect 483828 565528 485778 565584
rect 485834 565528 485839 565584
rect 483828 565526 485839 565528
rect 511796 565584 513439 565586
rect 511796 565528 513378 565584
rect 513434 565528 513439 565584
rect 511796 565526 513439 565528
rect 539948 565584 542419 565586
rect 539948 565528 542358 565584
rect 542414 565528 542419 565584
rect 539948 565526 542419 565528
rect 567916 565584 570019 565586
rect 567916 565528 569958 565584
rect 570014 565528 570019 565584
rect 567916 565526 570019 565528
rect 37917 565523 37983 565526
rect 66253 565523 66319 565526
rect 93853 565523 93919 565526
rect 121453 565523 121519 565526
rect 149053 565523 149119 565526
rect 178033 565523 178099 565526
rect 205633 565523 205699 565526
rect 233233 565523 233299 565526
rect 262213 565523 262279 565526
rect 289813 565523 289879 565526
rect 317413 565523 317479 565526
rect 345013 565523 345079 565526
rect 373993 565523 374059 565526
rect 401593 565523 401659 565526
rect 429193 565523 429259 565526
rect 458173 565523 458239 565526
rect 485773 565523 485839 565526
rect 513373 565523 513439 565526
rect 542353 565523 542419 565526
rect 569953 565523 570019 565526
rect 580257 564362 580323 564365
rect 583520 564362 584960 564452
rect 580257 564360 584960 564362
rect 580257 564304 580262 564360
rect 580318 564304 584960 564360
rect 580257 564302 584960 564304
rect 580257 564299 580323 564302
rect 583520 564212 584960 564302
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 13721 539338 13787 539341
rect 42701 539338 42767 539341
rect 70301 539338 70367 539341
rect 97901 539338 97967 539341
rect 126881 539338 126947 539341
rect 154481 539338 154547 539341
rect 182081 539338 182147 539341
rect 209681 539338 209747 539341
rect 238661 539338 238727 539341
rect 266261 539338 266327 539341
rect 293861 539338 293927 539341
rect 322841 539338 322907 539341
rect 350441 539338 350507 539341
rect 378041 539338 378107 539341
rect 405641 539338 405707 539341
rect 434621 539338 434687 539341
rect 462221 539338 462287 539341
rect 489821 539338 489887 539341
rect 518801 539338 518867 539341
rect 545757 539338 545823 539341
rect 13721 539336 16100 539338
rect 13721 539280 13726 539336
rect 13782 539280 16100 539336
rect 13721 539278 16100 539280
rect 42701 539336 44068 539338
rect 42701 539280 42706 539336
rect 42762 539280 44068 539336
rect 42701 539278 44068 539280
rect 70301 539336 72036 539338
rect 70301 539280 70306 539336
rect 70362 539280 72036 539336
rect 70301 539278 72036 539280
rect 97901 539336 100188 539338
rect 97901 539280 97906 539336
rect 97962 539280 100188 539336
rect 97901 539278 100188 539280
rect 126881 539336 128156 539338
rect 126881 539280 126886 539336
rect 126942 539280 128156 539336
rect 126881 539278 128156 539280
rect 154481 539336 156124 539338
rect 154481 539280 154486 539336
rect 154542 539280 156124 539336
rect 154481 539278 156124 539280
rect 182081 539336 184092 539338
rect 182081 539280 182086 539336
rect 182142 539280 184092 539336
rect 182081 539278 184092 539280
rect 209681 539336 212060 539338
rect 209681 539280 209686 539336
rect 209742 539280 212060 539336
rect 209681 539278 212060 539280
rect 238661 539336 240212 539338
rect 238661 539280 238666 539336
rect 238722 539280 240212 539336
rect 238661 539278 240212 539280
rect 266261 539336 268180 539338
rect 266261 539280 266266 539336
rect 266322 539280 268180 539336
rect 266261 539278 268180 539280
rect 293861 539336 296148 539338
rect 293861 539280 293866 539336
rect 293922 539280 296148 539336
rect 293861 539278 296148 539280
rect 322841 539336 324116 539338
rect 322841 539280 322846 539336
rect 322902 539280 324116 539336
rect 322841 539278 324116 539280
rect 350441 539336 352084 539338
rect 350441 539280 350446 539336
rect 350502 539280 352084 539336
rect 350441 539278 352084 539280
rect 378041 539336 380052 539338
rect 378041 539280 378046 539336
rect 378102 539280 380052 539336
rect 378041 539278 380052 539280
rect 405641 539336 408204 539338
rect 405641 539280 405646 539336
rect 405702 539280 408204 539336
rect 405641 539278 408204 539280
rect 434621 539336 436172 539338
rect 434621 539280 434626 539336
rect 434682 539280 436172 539336
rect 434621 539278 436172 539280
rect 462221 539336 464140 539338
rect 462221 539280 462226 539336
rect 462282 539280 464140 539336
rect 462221 539278 464140 539280
rect 489821 539336 492108 539338
rect 489821 539280 489826 539336
rect 489882 539280 492108 539336
rect 489821 539278 492108 539280
rect 518801 539336 520076 539338
rect 518801 539280 518806 539336
rect 518862 539280 520076 539336
rect 518801 539278 520076 539280
rect 545757 539336 548044 539338
rect 545757 539280 545762 539336
rect 545818 539280 548044 539336
rect 545757 539278 548044 539280
rect 13721 539275 13787 539278
rect 42701 539275 42767 539278
rect 70301 539275 70367 539278
rect 97901 539275 97967 539278
rect 126881 539275 126947 539278
rect 154481 539275 154547 539278
rect 182081 539275 182147 539278
rect 209681 539275 209747 539278
rect 238661 539275 238727 539278
rect 266261 539275 266327 539278
rect 293861 539275 293927 539278
rect 322841 539275 322907 539278
rect 350441 539275 350507 539278
rect 378041 539275 378107 539278
rect 405641 539275 405707 539278
rect 434621 539275 434687 539278
rect 462221 539275 462287 539278
rect 489821 539275 489887 539278
rect 518801 539275 518867 539278
rect 545757 539275 545823 539278
rect 37917 538658 37983 538661
rect 66253 538658 66319 538661
rect 93853 538658 93919 538661
rect 121453 538658 121519 538661
rect 149053 538658 149119 538661
rect 178033 538658 178099 538661
rect 205633 538658 205699 538661
rect 233233 538658 233299 538661
rect 262213 538658 262279 538661
rect 289813 538658 289879 538661
rect 317413 538658 317479 538661
rect 345013 538658 345079 538661
rect 373993 538658 374059 538661
rect 401593 538658 401659 538661
rect 429193 538658 429259 538661
rect 458173 538658 458239 538661
rect 485773 538658 485839 538661
rect 513373 538658 513439 538661
rect 542353 538658 542419 538661
rect 569953 538658 570019 538661
rect 35788 538656 37983 538658
rect 35788 538600 37922 538656
rect 37978 538600 37983 538656
rect 35788 538598 37983 538600
rect 63940 538656 66319 538658
rect 63940 538600 66258 538656
rect 66314 538600 66319 538656
rect 63940 538598 66319 538600
rect 91908 538656 93919 538658
rect 91908 538600 93858 538656
rect 93914 538600 93919 538656
rect 91908 538598 93919 538600
rect 119876 538656 121519 538658
rect 119876 538600 121458 538656
rect 121514 538600 121519 538656
rect 119876 538598 121519 538600
rect 147844 538656 149119 538658
rect 147844 538600 149058 538656
rect 149114 538600 149119 538656
rect 147844 538598 149119 538600
rect 175812 538656 178099 538658
rect 175812 538600 178038 538656
rect 178094 538600 178099 538656
rect 175812 538598 178099 538600
rect 203964 538656 205699 538658
rect 203964 538600 205638 538656
rect 205694 538600 205699 538656
rect 203964 538598 205699 538600
rect 231932 538656 233299 538658
rect 231932 538600 233238 538656
rect 233294 538600 233299 538656
rect 231932 538598 233299 538600
rect 259900 538656 262279 538658
rect 259900 538600 262218 538656
rect 262274 538600 262279 538656
rect 259900 538598 262279 538600
rect 287868 538656 289879 538658
rect 287868 538600 289818 538656
rect 289874 538600 289879 538656
rect 287868 538598 289879 538600
rect 315836 538656 317479 538658
rect 315836 538600 317418 538656
rect 317474 538600 317479 538656
rect 315836 538598 317479 538600
rect 343804 538656 345079 538658
rect 343804 538600 345018 538656
rect 345074 538600 345079 538656
rect 343804 538598 345079 538600
rect 371956 538656 374059 538658
rect 371956 538600 373998 538656
rect 374054 538600 374059 538656
rect 371956 538598 374059 538600
rect 399924 538656 401659 538658
rect 399924 538600 401598 538656
rect 401654 538600 401659 538656
rect 399924 538598 401659 538600
rect 427892 538656 429259 538658
rect 427892 538600 429198 538656
rect 429254 538600 429259 538656
rect 427892 538598 429259 538600
rect 455860 538656 458239 538658
rect 455860 538600 458178 538656
rect 458234 538600 458239 538656
rect 455860 538598 458239 538600
rect 483828 538656 485839 538658
rect 483828 538600 485778 538656
rect 485834 538600 485839 538656
rect 483828 538598 485839 538600
rect 511796 538656 513439 538658
rect 511796 538600 513378 538656
rect 513434 538600 513439 538656
rect 511796 538598 513439 538600
rect 539948 538656 542419 538658
rect 539948 538600 542358 538656
rect 542414 538600 542419 538656
rect 539948 538598 542419 538600
rect 567916 538656 570019 538658
rect 567916 538600 569958 538656
rect 570014 538600 570019 538656
rect 567916 538598 570019 538600
rect 37917 538595 37983 538598
rect 66253 538595 66319 538598
rect 93853 538595 93919 538598
rect 121453 538595 121519 538598
rect 149053 538595 149119 538598
rect 178033 538595 178099 538598
rect 205633 538595 205699 538598
rect 233233 538595 233299 538598
rect 262213 538595 262279 538598
rect 289813 538595 289879 538598
rect 317413 538595 317479 538598
rect 345013 538595 345079 538598
rect 373993 538595 374059 538598
rect 401593 538595 401659 538598
rect 429193 538595 429259 538598
rect 458173 538595 458239 538598
rect 485773 538595 485839 538598
rect 513373 538595 513439 538598
rect 542353 538595 542419 538598
rect 569953 538595 570019 538598
rect 583520 537692 584960 537932
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 407849 512818 407915 512821
rect 407849 512816 408234 512818
rect 407849 512760 407854 512816
rect 407910 512760 408234 512816
rect 407849 512758 408234 512760
rect 407849 512755 407915 512758
rect 13721 512274 13787 512277
rect 42701 512274 42767 512277
rect 70301 512274 70367 512277
rect 97901 512274 97967 512277
rect 126881 512274 126947 512277
rect 154481 512274 154547 512277
rect 182081 512274 182147 512277
rect 209681 512274 209747 512277
rect 238661 512274 238727 512277
rect 266261 512274 266327 512277
rect 293861 512274 293927 512277
rect 322841 512274 322907 512277
rect 350441 512274 350507 512277
rect 378041 512274 378107 512277
rect 13721 512272 16100 512274
rect 13721 512216 13726 512272
rect 13782 512216 16100 512272
rect 13721 512214 16100 512216
rect 42701 512272 44068 512274
rect 42701 512216 42706 512272
rect 42762 512216 44068 512272
rect 42701 512214 44068 512216
rect 70301 512272 72036 512274
rect 70301 512216 70306 512272
rect 70362 512216 72036 512272
rect 70301 512214 72036 512216
rect 97901 512272 100188 512274
rect 97901 512216 97906 512272
rect 97962 512216 100188 512272
rect 97901 512214 100188 512216
rect 126881 512272 128156 512274
rect 126881 512216 126886 512272
rect 126942 512216 128156 512272
rect 126881 512214 128156 512216
rect 154481 512272 156124 512274
rect 154481 512216 154486 512272
rect 154542 512216 156124 512272
rect 154481 512214 156124 512216
rect 182081 512272 184092 512274
rect 182081 512216 182086 512272
rect 182142 512216 184092 512272
rect 182081 512214 184092 512216
rect 209681 512272 212060 512274
rect 209681 512216 209686 512272
rect 209742 512216 212060 512272
rect 209681 512214 212060 512216
rect 238661 512272 240212 512274
rect 238661 512216 238666 512272
rect 238722 512216 240212 512272
rect 238661 512214 240212 512216
rect 266261 512272 268180 512274
rect 266261 512216 266266 512272
rect 266322 512216 268180 512272
rect 266261 512214 268180 512216
rect 293861 512272 296148 512274
rect 293861 512216 293866 512272
rect 293922 512216 296148 512272
rect 293861 512214 296148 512216
rect 322841 512272 324116 512274
rect 322841 512216 322846 512272
rect 322902 512216 324116 512272
rect 322841 512214 324116 512216
rect 350441 512272 352084 512274
rect 350441 512216 350446 512272
rect 350502 512216 352084 512272
rect 350441 512214 352084 512216
rect 378041 512272 380052 512274
rect 378041 512216 378046 512272
rect 378102 512216 380052 512272
rect 408174 512244 408234 512758
rect 434621 512274 434687 512277
rect 462221 512274 462287 512277
rect 489821 512274 489887 512277
rect 518801 512274 518867 512277
rect 545757 512274 545823 512277
rect 434621 512272 436172 512274
rect 378041 512214 380052 512216
rect 434621 512216 434626 512272
rect 434682 512216 436172 512272
rect 434621 512214 436172 512216
rect 462221 512272 464140 512274
rect 462221 512216 462226 512272
rect 462282 512216 464140 512272
rect 462221 512214 464140 512216
rect 489821 512272 492108 512274
rect 489821 512216 489826 512272
rect 489882 512216 492108 512272
rect 489821 512214 492108 512216
rect 518801 512272 520076 512274
rect 518801 512216 518806 512272
rect 518862 512216 520076 512272
rect 518801 512214 520076 512216
rect 545757 512272 548044 512274
rect 545757 512216 545762 512272
rect 545818 512216 548044 512272
rect 545757 512214 548044 512216
rect 13721 512211 13787 512214
rect 42701 512211 42767 512214
rect 70301 512211 70367 512214
rect 97901 512211 97967 512214
rect 126881 512211 126947 512214
rect 154481 512211 154547 512214
rect 182081 512211 182147 512214
rect 209681 512211 209747 512214
rect 238661 512211 238727 512214
rect 266261 512211 266327 512214
rect 293861 512211 293927 512214
rect 322841 512211 322907 512214
rect 350441 512211 350507 512214
rect 378041 512211 378107 512214
rect 434621 512211 434687 512214
rect 462221 512211 462287 512214
rect 489821 512211 489887 512214
rect 518801 512211 518867 512214
rect 545757 512211 545823 512214
rect 37917 511594 37983 511597
rect 66253 511594 66319 511597
rect 93853 511594 93919 511597
rect 121453 511594 121519 511597
rect 149053 511594 149119 511597
rect 178033 511594 178099 511597
rect 205633 511594 205699 511597
rect 233233 511594 233299 511597
rect 262213 511594 262279 511597
rect 289813 511594 289879 511597
rect 317413 511594 317479 511597
rect 345013 511594 345079 511597
rect 373993 511594 374059 511597
rect 401593 511594 401659 511597
rect 429193 511594 429259 511597
rect 458173 511594 458239 511597
rect 485773 511594 485839 511597
rect 513373 511594 513439 511597
rect 569953 511594 570019 511597
rect 35788 511592 37983 511594
rect 35788 511536 37922 511592
rect 37978 511536 37983 511592
rect 35788 511534 37983 511536
rect 63940 511592 66319 511594
rect 63940 511536 66258 511592
rect 66314 511536 66319 511592
rect 63940 511534 66319 511536
rect 91908 511592 93919 511594
rect 91908 511536 93858 511592
rect 93914 511536 93919 511592
rect 91908 511534 93919 511536
rect 119876 511592 121519 511594
rect 119876 511536 121458 511592
rect 121514 511536 121519 511592
rect 119876 511534 121519 511536
rect 147844 511592 149119 511594
rect 147844 511536 149058 511592
rect 149114 511536 149119 511592
rect 147844 511534 149119 511536
rect 175812 511592 178099 511594
rect 175812 511536 178038 511592
rect 178094 511536 178099 511592
rect 175812 511534 178099 511536
rect 203964 511592 205699 511594
rect 203964 511536 205638 511592
rect 205694 511536 205699 511592
rect 203964 511534 205699 511536
rect 231932 511592 233299 511594
rect 231932 511536 233238 511592
rect 233294 511536 233299 511592
rect 231932 511534 233299 511536
rect 259900 511592 262279 511594
rect 259900 511536 262218 511592
rect 262274 511536 262279 511592
rect 259900 511534 262279 511536
rect 287868 511592 289879 511594
rect 287868 511536 289818 511592
rect 289874 511536 289879 511592
rect 287868 511534 289879 511536
rect 315836 511592 317479 511594
rect 315836 511536 317418 511592
rect 317474 511536 317479 511592
rect 315836 511534 317479 511536
rect 343804 511592 345079 511594
rect 343804 511536 345018 511592
rect 345074 511536 345079 511592
rect 343804 511534 345079 511536
rect 371956 511592 374059 511594
rect 371956 511536 373998 511592
rect 374054 511536 374059 511592
rect 371956 511534 374059 511536
rect 399924 511592 401659 511594
rect 399924 511536 401598 511592
rect 401654 511536 401659 511592
rect 399924 511534 401659 511536
rect 427892 511592 429259 511594
rect 427892 511536 429198 511592
rect 429254 511536 429259 511592
rect 427892 511534 429259 511536
rect 455860 511592 458239 511594
rect 455860 511536 458178 511592
rect 458234 511536 458239 511592
rect 455860 511534 458239 511536
rect 483828 511592 485839 511594
rect 483828 511536 485778 511592
rect 485834 511536 485839 511592
rect 483828 511534 485839 511536
rect 511796 511592 513439 511594
rect 511796 511536 513378 511592
rect 513434 511536 513439 511592
rect 567916 511592 570019 511594
rect 511796 511534 513439 511536
rect 37917 511531 37983 511534
rect 66253 511531 66319 511534
rect 93853 511531 93919 511534
rect 121453 511531 121519 511534
rect 149053 511531 149119 511534
rect 178033 511531 178099 511534
rect 205633 511531 205699 511534
rect 233233 511531 233299 511534
rect 262213 511531 262279 511534
rect 289813 511531 289879 511534
rect 317413 511531 317479 511534
rect 345013 511531 345079 511534
rect 373993 511531 374059 511534
rect 401593 511531 401659 511534
rect 429193 511531 429259 511534
rect 458173 511531 458239 511534
rect 485773 511531 485839 511534
rect 513373 511531 513439 511534
rect 539918 511050 539978 511564
rect 567916 511536 569958 511592
rect 570014 511536 570019 511592
rect 567916 511534 570019 511536
rect 569953 511531 570019 511534
rect 583520 511172 584960 511412
rect 540881 511050 540947 511053
rect 539918 511048 540947 511050
rect 539918 510992 540886 511048
rect 540942 510992 540947 511048
rect 539918 510990 540947 510992
rect 540881 510987 540947 510990
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 13721 485346 13787 485349
rect 42701 485346 42767 485349
rect 97901 485346 97967 485349
rect 126881 485346 126947 485349
rect 154481 485346 154547 485349
rect 182081 485346 182147 485349
rect 209681 485346 209747 485349
rect 238661 485346 238727 485349
rect 266261 485346 266327 485349
rect 293861 485346 293927 485349
rect 322841 485346 322907 485349
rect 350441 485346 350507 485349
rect 378041 485346 378107 485349
rect 405641 485346 405707 485349
rect 434621 485346 434687 485349
rect 462221 485346 462287 485349
rect 489821 485346 489887 485349
rect 518801 485346 518867 485349
rect 545757 485346 545823 485349
rect 13721 485344 16100 485346
rect 13721 485288 13726 485344
rect 13782 485288 16100 485344
rect 13721 485286 16100 485288
rect 42701 485344 44068 485346
rect 42701 485288 42706 485344
rect 42762 485288 44068 485344
rect 97901 485344 100188 485346
rect 42701 485286 44068 485288
rect 13721 485283 13787 485286
rect 42701 485283 42767 485286
rect 70301 484802 70367 484805
rect 72006 484802 72066 485316
rect 97901 485288 97906 485344
rect 97962 485288 100188 485344
rect 97901 485286 100188 485288
rect 126881 485344 128156 485346
rect 126881 485288 126886 485344
rect 126942 485288 128156 485344
rect 126881 485286 128156 485288
rect 154481 485344 156124 485346
rect 154481 485288 154486 485344
rect 154542 485288 156124 485344
rect 154481 485286 156124 485288
rect 182081 485344 184092 485346
rect 182081 485288 182086 485344
rect 182142 485288 184092 485344
rect 182081 485286 184092 485288
rect 209681 485344 212060 485346
rect 209681 485288 209686 485344
rect 209742 485288 212060 485344
rect 209681 485286 212060 485288
rect 238661 485344 240212 485346
rect 238661 485288 238666 485344
rect 238722 485288 240212 485344
rect 238661 485286 240212 485288
rect 266261 485344 268180 485346
rect 266261 485288 266266 485344
rect 266322 485288 268180 485344
rect 266261 485286 268180 485288
rect 293861 485344 296148 485346
rect 293861 485288 293866 485344
rect 293922 485288 296148 485344
rect 293861 485286 296148 485288
rect 322841 485344 324116 485346
rect 322841 485288 322846 485344
rect 322902 485288 324116 485344
rect 322841 485286 324116 485288
rect 350441 485344 352084 485346
rect 350441 485288 350446 485344
rect 350502 485288 352084 485344
rect 350441 485286 352084 485288
rect 378041 485344 380052 485346
rect 378041 485288 378046 485344
rect 378102 485288 380052 485344
rect 378041 485286 380052 485288
rect 405641 485344 408204 485346
rect 405641 485288 405646 485344
rect 405702 485288 408204 485344
rect 405641 485286 408204 485288
rect 434621 485344 436172 485346
rect 434621 485288 434626 485344
rect 434682 485288 436172 485344
rect 434621 485286 436172 485288
rect 462221 485344 464140 485346
rect 462221 485288 462226 485344
rect 462282 485288 464140 485344
rect 462221 485286 464140 485288
rect 489821 485344 492108 485346
rect 489821 485288 489826 485344
rect 489882 485288 492108 485344
rect 489821 485286 492108 485288
rect 518801 485344 520076 485346
rect 518801 485288 518806 485344
rect 518862 485288 520076 485344
rect 518801 485286 520076 485288
rect 545757 485344 548044 485346
rect 545757 485288 545762 485344
rect 545818 485288 548044 485344
rect 545757 485286 548044 485288
rect 97901 485283 97967 485286
rect 126881 485283 126947 485286
rect 154481 485283 154547 485286
rect 182081 485283 182147 485286
rect 209681 485283 209747 485286
rect 238661 485283 238727 485286
rect 266261 485283 266327 485286
rect 293861 485283 293927 485286
rect 322841 485283 322907 485286
rect 350441 485283 350507 485286
rect 378041 485283 378107 485286
rect 405641 485283 405707 485286
rect 434621 485283 434687 485286
rect 462221 485283 462287 485286
rect 489821 485283 489887 485286
rect 518801 485283 518867 485286
rect 545757 485283 545823 485286
rect 70301 484800 72066 484802
rect 70301 484744 70306 484800
rect 70362 484744 72066 484800
rect 70301 484742 72066 484744
rect 70301 484739 70367 484742
rect 37917 484666 37983 484669
rect 66253 484666 66319 484669
rect 93853 484666 93919 484669
rect 121453 484666 121519 484669
rect 149053 484666 149119 484669
rect 178033 484666 178099 484669
rect 233233 484666 233299 484669
rect 262213 484666 262279 484669
rect 289813 484666 289879 484669
rect 317413 484666 317479 484669
rect 345013 484666 345079 484669
rect 373993 484666 374059 484669
rect 401593 484666 401659 484669
rect 429193 484666 429259 484669
rect 458173 484666 458239 484669
rect 485773 484666 485839 484669
rect 513373 484666 513439 484669
rect 542353 484666 542419 484669
rect 569953 484666 570019 484669
rect 35788 484664 37983 484666
rect 35788 484608 37922 484664
rect 37978 484608 37983 484664
rect 35788 484606 37983 484608
rect 63940 484664 66319 484666
rect 63940 484608 66258 484664
rect 66314 484608 66319 484664
rect 63940 484606 66319 484608
rect 91908 484664 93919 484666
rect 91908 484608 93858 484664
rect 93914 484608 93919 484664
rect 91908 484606 93919 484608
rect 119876 484664 121519 484666
rect 119876 484608 121458 484664
rect 121514 484608 121519 484664
rect 119876 484606 121519 484608
rect 147844 484664 149119 484666
rect 147844 484608 149058 484664
rect 149114 484608 149119 484664
rect 147844 484606 149119 484608
rect 175812 484664 178099 484666
rect 175812 484608 178038 484664
rect 178094 484608 178099 484664
rect 231932 484664 233299 484666
rect 175812 484606 178099 484608
rect 37917 484603 37983 484606
rect 66253 484603 66319 484606
rect 93853 484603 93919 484606
rect 121453 484603 121519 484606
rect 149053 484603 149119 484606
rect 178033 484603 178099 484606
rect 203934 484530 203994 484636
rect 231932 484608 233238 484664
rect 233294 484608 233299 484664
rect 231932 484606 233299 484608
rect 259900 484664 262279 484666
rect 259900 484608 262218 484664
rect 262274 484608 262279 484664
rect 259900 484606 262279 484608
rect 287868 484664 289879 484666
rect 287868 484608 289818 484664
rect 289874 484608 289879 484664
rect 287868 484606 289879 484608
rect 315836 484664 317479 484666
rect 315836 484608 317418 484664
rect 317474 484608 317479 484664
rect 315836 484606 317479 484608
rect 343804 484664 345079 484666
rect 343804 484608 345018 484664
rect 345074 484608 345079 484664
rect 343804 484606 345079 484608
rect 371956 484664 374059 484666
rect 371956 484608 373998 484664
rect 374054 484608 374059 484664
rect 371956 484606 374059 484608
rect 399924 484664 401659 484666
rect 399924 484608 401598 484664
rect 401654 484608 401659 484664
rect 399924 484606 401659 484608
rect 427892 484664 429259 484666
rect 427892 484608 429198 484664
rect 429254 484608 429259 484664
rect 427892 484606 429259 484608
rect 455860 484664 458239 484666
rect 455860 484608 458178 484664
rect 458234 484608 458239 484664
rect 455860 484606 458239 484608
rect 483828 484664 485839 484666
rect 483828 484608 485778 484664
rect 485834 484608 485839 484664
rect 483828 484606 485839 484608
rect 511796 484664 513439 484666
rect 511796 484608 513378 484664
rect 513434 484608 513439 484664
rect 511796 484606 513439 484608
rect 539948 484664 542419 484666
rect 539948 484608 542358 484664
rect 542414 484608 542419 484664
rect 539948 484606 542419 484608
rect 567916 484664 570019 484666
rect 567916 484608 569958 484664
rect 570014 484608 570019 484664
rect 567916 484606 570019 484608
rect 233233 484603 233299 484606
rect 262213 484603 262279 484606
rect 289813 484603 289879 484606
rect 317413 484603 317479 484606
rect 345013 484603 345079 484606
rect 373993 484603 374059 484606
rect 401593 484603 401659 484606
rect 429193 484603 429259 484606
rect 458173 484603 458239 484606
rect 485773 484603 485839 484606
rect 513373 484603 513439 484606
rect 542353 484603 542419 484606
rect 569953 484603 570019 484606
rect 205633 484530 205699 484533
rect 203934 484528 205699 484530
rect 203934 484472 205638 484528
rect 205694 484472 205699 484528
rect 583520 484516 584960 484756
rect 203934 484470 205699 484472
rect 205633 484467 205699 484470
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 13721 458282 13787 458285
rect 42701 458282 42767 458285
rect 70301 458282 70367 458285
rect 97901 458282 97967 458285
rect 126881 458282 126947 458285
rect 154481 458282 154547 458285
rect 182081 458282 182147 458285
rect 209681 458282 209747 458285
rect 238661 458282 238727 458285
rect 266261 458282 266327 458285
rect 293861 458282 293927 458285
rect 322841 458282 322907 458285
rect 350441 458282 350507 458285
rect 378041 458282 378107 458285
rect 405641 458282 405707 458285
rect 434621 458282 434687 458285
rect 462221 458282 462287 458285
rect 489821 458282 489887 458285
rect 518801 458282 518867 458285
rect 545757 458282 545823 458285
rect 13721 458280 16100 458282
rect 13721 458224 13726 458280
rect 13782 458224 16100 458280
rect 13721 458222 16100 458224
rect 42701 458280 44068 458282
rect 42701 458224 42706 458280
rect 42762 458224 44068 458280
rect 42701 458222 44068 458224
rect 70301 458280 72036 458282
rect 70301 458224 70306 458280
rect 70362 458224 72036 458280
rect 70301 458222 72036 458224
rect 97901 458280 100188 458282
rect 97901 458224 97906 458280
rect 97962 458224 100188 458280
rect 97901 458222 100188 458224
rect 126881 458280 128156 458282
rect 126881 458224 126886 458280
rect 126942 458224 128156 458280
rect 126881 458222 128156 458224
rect 154481 458280 156124 458282
rect 154481 458224 154486 458280
rect 154542 458224 156124 458280
rect 154481 458222 156124 458224
rect 182081 458280 184092 458282
rect 182081 458224 182086 458280
rect 182142 458224 184092 458280
rect 182081 458222 184092 458224
rect 209681 458280 212060 458282
rect 209681 458224 209686 458280
rect 209742 458224 212060 458280
rect 209681 458222 212060 458224
rect 238661 458280 240212 458282
rect 238661 458224 238666 458280
rect 238722 458224 240212 458280
rect 238661 458222 240212 458224
rect 266261 458280 268180 458282
rect 266261 458224 266266 458280
rect 266322 458224 268180 458280
rect 266261 458222 268180 458224
rect 293861 458280 296148 458282
rect 293861 458224 293866 458280
rect 293922 458224 296148 458280
rect 293861 458222 296148 458224
rect 322841 458280 324116 458282
rect 322841 458224 322846 458280
rect 322902 458224 324116 458280
rect 322841 458222 324116 458224
rect 350441 458280 352084 458282
rect 350441 458224 350446 458280
rect 350502 458224 352084 458280
rect 350441 458222 352084 458224
rect 378041 458280 380052 458282
rect 378041 458224 378046 458280
rect 378102 458224 380052 458280
rect 378041 458222 380052 458224
rect 405641 458280 408204 458282
rect 405641 458224 405646 458280
rect 405702 458224 408204 458280
rect 405641 458222 408204 458224
rect 434621 458280 436172 458282
rect 434621 458224 434626 458280
rect 434682 458224 436172 458280
rect 434621 458222 436172 458224
rect 462221 458280 464140 458282
rect 462221 458224 462226 458280
rect 462282 458224 464140 458280
rect 462221 458222 464140 458224
rect 489821 458280 492108 458282
rect 489821 458224 489826 458280
rect 489882 458224 492108 458280
rect 489821 458222 492108 458224
rect 518801 458280 520076 458282
rect 518801 458224 518806 458280
rect 518862 458224 520076 458280
rect 518801 458222 520076 458224
rect 545757 458280 548044 458282
rect 545757 458224 545762 458280
rect 545818 458224 548044 458280
rect 545757 458222 548044 458224
rect 13721 458219 13787 458222
rect 42701 458219 42767 458222
rect 70301 458219 70367 458222
rect 97901 458219 97967 458222
rect 126881 458219 126947 458222
rect 154481 458219 154547 458222
rect 182081 458219 182147 458222
rect 209681 458219 209747 458222
rect 238661 458219 238727 458222
rect 266261 458219 266327 458222
rect 293861 458219 293927 458222
rect 322841 458219 322907 458222
rect 350441 458219 350507 458222
rect 378041 458219 378107 458222
rect 405641 458219 405707 458222
rect 434621 458219 434687 458222
rect 462221 458219 462287 458222
rect 489821 458219 489887 458222
rect 518801 458219 518867 458222
rect 545757 458219 545823 458222
rect 583520 457996 584960 458236
rect 37917 457602 37983 457605
rect 66253 457602 66319 457605
rect 93853 457602 93919 457605
rect 121453 457602 121519 457605
rect 149053 457602 149119 457605
rect 178033 457602 178099 457605
rect 205633 457602 205699 457605
rect 233233 457602 233299 457605
rect 262213 457602 262279 457605
rect 289813 457602 289879 457605
rect 317413 457602 317479 457605
rect 345013 457602 345079 457605
rect 373993 457602 374059 457605
rect 401593 457602 401659 457605
rect 429193 457602 429259 457605
rect 458173 457602 458239 457605
rect 485773 457602 485839 457605
rect 513373 457602 513439 457605
rect 542353 457602 542419 457605
rect 569953 457602 570019 457605
rect 35788 457600 37983 457602
rect 35788 457544 37922 457600
rect 37978 457544 37983 457600
rect 35788 457542 37983 457544
rect 63940 457600 66319 457602
rect 63940 457544 66258 457600
rect 66314 457544 66319 457600
rect 63940 457542 66319 457544
rect 91908 457600 93919 457602
rect 91908 457544 93858 457600
rect 93914 457544 93919 457600
rect 91908 457542 93919 457544
rect 119876 457600 121519 457602
rect 119876 457544 121458 457600
rect 121514 457544 121519 457600
rect 119876 457542 121519 457544
rect 147844 457600 149119 457602
rect 147844 457544 149058 457600
rect 149114 457544 149119 457600
rect 147844 457542 149119 457544
rect 175812 457600 178099 457602
rect 175812 457544 178038 457600
rect 178094 457544 178099 457600
rect 175812 457542 178099 457544
rect 203964 457600 205699 457602
rect 203964 457544 205638 457600
rect 205694 457544 205699 457600
rect 203964 457542 205699 457544
rect 231932 457600 233299 457602
rect 231932 457544 233238 457600
rect 233294 457544 233299 457600
rect 231932 457542 233299 457544
rect 259900 457600 262279 457602
rect 259900 457544 262218 457600
rect 262274 457544 262279 457600
rect 259900 457542 262279 457544
rect 287868 457600 289879 457602
rect 287868 457544 289818 457600
rect 289874 457544 289879 457600
rect 287868 457542 289879 457544
rect 315836 457600 317479 457602
rect 315836 457544 317418 457600
rect 317474 457544 317479 457600
rect 315836 457542 317479 457544
rect 343804 457600 345079 457602
rect 343804 457544 345018 457600
rect 345074 457544 345079 457600
rect 343804 457542 345079 457544
rect 371956 457600 374059 457602
rect 371956 457544 373998 457600
rect 374054 457544 374059 457600
rect 371956 457542 374059 457544
rect 399924 457600 401659 457602
rect 399924 457544 401598 457600
rect 401654 457544 401659 457600
rect 399924 457542 401659 457544
rect 427892 457600 429259 457602
rect 427892 457544 429198 457600
rect 429254 457544 429259 457600
rect 427892 457542 429259 457544
rect 455860 457600 458239 457602
rect 455860 457544 458178 457600
rect 458234 457544 458239 457600
rect 455860 457542 458239 457544
rect 483828 457600 485839 457602
rect 483828 457544 485778 457600
rect 485834 457544 485839 457600
rect 483828 457542 485839 457544
rect 511796 457600 513439 457602
rect 511796 457544 513378 457600
rect 513434 457544 513439 457600
rect 511796 457542 513439 457544
rect 539948 457600 542419 457602
rect 539948 457544 542358 457600
rect 542414 457544 542419 457600
rect 539948 457542 542419 457544
rect 567916 457600 570019 457602
rect 567916 457544 569958 457600
rect 570014 457544 570019 457600
rect 567916 457542 570019 457544
rect 37917 457539 37983 457542
rect 66253 457539 66319 457542
rect 93853 457539 93919 457542
rect 121453 457539 121519 457542
rect 149053 457539 149119 457542
rect 178033 457539 178099 457542
rect 205633 457539 205699 457542
rect 233233 457539 233299 457542
rect 262213 457539 262279 457542
rect 289813 457539 289879 457542
rect 317413 457539 317479 457542
rect 345013 457539 345079 457542
rect 373993 457539 374059 457542
rect 401593 457539 401659 457542
rect 429193 457539 429259 457542
rect 458173 457539 458239 457542
rect 485773 457539 485839 457542
rect 513373 457539 513439 457542
rect 542353 457539 542419 457542
rect 569953 457539 570019 457542
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 545757 431898 545823 431901
rect 545757 431896 548074 431898
rect 545757 431840 545762 431896
rect 545818 431840 548074 431896
rect 545757 431838 548074 431840
rect 545757 431835 545823 431838
rect 13721 431354 13787 431357
rect 42701 431354 42767 431357
rect 97901 431354 97967 431357
rect 126881 431354 126947 431357
rect 154481 431354 154547 431357
rect 182081 431354 182147 431357
rect 209681 431354 209747 431357
rect 238661 431354 238727 431357
rect 266261 431354 266327 431357
rect 293861 431354 293927 431357
rect 322841 431354 322907 431357
rect 350441 431354 350507 431357
rect 378041 431354 378107 431357
rect 405641 431354 405707 431357
rect 434621 431354 434687 431357
rect 462221 431354 462287 431357
rect 489821 431354 489887 431357
rect 518801 431354 518867 431357
rect 13721 431352 16100 431354
rect 13721 431296 13726 431352
rect 13782 431296 16100 431352
rect 13721 431294 16100 431296
rect 42701 431352 44068 431354
rect 42701 431296 42706 431352
rect 42762 431296 44068 431352
rect 97901 431352 100188 431354
rect 42701 431294 44068 431296
rect 13721 431291 13787 431294
rect 42701 431291 42767 431294
rect 70301 430810 70367 430813
rect 72006 430810 72066 431324
rect 97901 431296 97906 431352
rect 97962 431296 100188 431352
rect 97901 431294 100188 431296
rect 126881 431352 128156 431354
rect 126881 431296 126886 431352
rect 126942 431296 128156 431352
rect 126881 431294 128156 431296
rect 154481 431352 156124 431354
rect 154481 431296 154486 431352
rect 154542 431296 156124 431352
rect 154481 431294 156124 431296
rect 182081 431352 184092 431354
rect 182081 431296 182086 431352
rect 182142 431296 184092 431352
rect 182081 431294 184092 431296
rect 209681 431352 212060 431354
rect 209681 431296 209686 431352
rect 209742 431296 212060 431352
rect 209681 431294 212060 431296
rect 238661 431352 240212 431354
rect 238661 431296 238666 431352
rect 238722 431296 240212 431352
rect 238661 431294 240212 431296
rect 266261 431352 268180 431354
rect 266261 431296 266266 431352
rect 266322 431296 268180 431352
rect 266261 431294 268180 431296
rect 293861 431352 296148 431354
rect 293861 431296 293866 431352
rect 293922 431296 296148 431352
rect 293861 431294 296148 431296
rect 322841 431352 324116 431354
rect 322841 431296 322846 431352
rect 322902 431296 324116 431352
rect 322841 431294 324116 431296
rect 350441 431352 352084 431354
rect 350441 431296 350446 431352
rect 350502 431296 352084 431352
rect 350441 431294 352084 431296
rect 378041 431352 380052 431354
rect 378041 431296 378046 431352
rect 378102 431296 380052 431352
rect 378041 431294 380052 431296
rect 405641 431352 408204 431354
rect 405641 431296 405646 431352
rect 405702 431296 408204 431352
rect 405641 431294 408204 431296
rect 434621 431352 436172 431354
rect 434621 431296 434626 431352
rect 434682 431296 436172 431352
rect 434621 431294 436172 431296
rect 462221 431352 464140 431354
rect 462221 431296 462226 431352
rect 462282 431296 464140 431352
rect 462221 431294 464140 431296
rect 489821 431352 492108 431354
rect 489821 431296 489826 431352
rect 489882 431296 492108 431352
rect 489821 431294 492108 431296
rect 518801 431352 520076 431354
rect 518801 431296 518806 431352
rect 518862 431296 520076 431352
rect 548014 431324 548074 431838
rect 583520 431476 584960 431716
rect 518801 431294 520076 431296
rect 97901 431291 97967 431294
rect 126881 431291 126947 431294
rect 154481 431291 154547 431294
rect 182081 431291 182147 431294
rect 209681 431291 209747 431294
rect 238661 431291 238727 431294
rect 266261 431291 266327 431294
rect 293861 431291 293927 431294
rect 322841 431291 322907 431294
rect 350441 431291 350507 431294
rect 378041 431291 378107 431294
rect 405641 431291 405707 431294
rect 434621 431291 434687 431294
rect 462221 431291 462287 431294
rect 489821 431291 489887 431294
rect 518801 431291 518867 431294
rect 205633 431218 205699 431221
rect 70301 430808 72066 430810
rect 70301 430752 70306 430808
rect 70362 430752 72066 430808
rect 70301 430750 72066 430752
rect 203934 431216 205699 431218
rect 203934 431160 205638 431216
rect 205694 431160 205699 431216
rect 203934 431158 205699 431160
rect 70301 430747 70367 430750
rect 37917 430674 37983 430677
rect 66253 430674 66319 430677
rect 93853 430674 93919 430677
rect 121453 430674 121519 430677
rect 149053 430674 149119 430677
rect 178033 430674 178099 430677
rect 35788 430672 37983 430674
rect 35788 430616 37922 430672
rect 37978 430616 37983 430672
rect 35788 430614 37983 430616
rect 63940 430672 66319 430674
rect 63940 430616 66258 430672
rect 66314 430616 66319 430672
rect 63940 430614 66319 430616
rect 91908 430672 93919 430674
rect 91908 430616 93858 430672
rect 93914 430616 93919 430672
rect 91908 430614 93919 430616
rect 119876 430672 121519 430674
rect 119876 430616 121458 430672
rect 121514 430616 121519 430672
rect 119876 430614 121519 430616
rect 147844 430672 149119 430674
rect 147844 430616 149058 430672
rect 149114 430616 149119 430672
rect 147844 430614 149119 430616
rect 175812 430672 178099 430674
rect 175812 430616 178038 430672
rect 178094 430616 178099 430672
rect 203934 430644 203994 431158
rect 205633 431155 205699 431158
rect 373993 430810 374059 430813
rect 371926 430808 374059 430810
rect 371926 430752 373998 430808
rect 374054 430752 374059 430808
rect 371926 430750 374059 430752
rect 233233 430674 233299 430677
rect 262213 430674 262279 430677
rect 289813 430674 289879 430677
rect 317413 430674 317479 430677
rect 345013 430674 345079 430677
rect 231932 430672 233299 430674
rect 175812 430614 178099 430616
rect 231932 430616 233238 430672
rect 233294 430616 233299 430672
rect 231932 430614 233299 430616
rect 259900 430672 262279 430674
rect 259900 430616 262218 430672
rect 262274 430616 262279 430672
rect 259900 430614 262279 430616
rect 287868 430672 289879 430674
rect 287868 430616 289818 430672
rect 289874 430616 289879 430672
rect 287868 430614 289879 430616
rect 315836 430672 317479 430674
rect 315836 430616 317418 430672
rect 317474 430616 317479 430672
rect 315836 430614 317479 430616
rect 343804 430672 345079 430674
rect 343804 430616 345018 430672
rect 345074 430616 345079 430672
rect 371926 430644 371986 430750
rect 373993 430747 374059 430750
rect 401593 430674 401659 430677
rect 429193 430674 429259 430677
rect 458173 430674 458239 430677
rect 485773 430674 485839 430677
rect 513373 430674 513439 430677
rect 542353 430674 542419 430677
rect 569953 430674 570019 430677
rect 399924 430672 401659 430674
rect 343804 430614 345079 430616
rect 399924 430616 401598 430672
rect 401654 430616 401659 430672
rect 399924 430614 401659 430616
rect 427892 430672 429259 430674
rect 427892 430616 429198 430672
rect 429254 430616 429259 430672
rect 427892 430614 429259 430616
rect 455860 430672 458239 430674
rect 455860 430616 458178 430672
rect 458234 430616 458239 430672
rect 455860 430614 458239 430616
rect 483828 430672 485839 430674
rect 483828 430616 485778 430672
rect 485834 430616 485839 430672
rect 483828 430614 485839 430616
rect 511796 430672 513439 430674
rect 511796 430616 513378 430672
rect 513434 430616 513439 430672
rect 511796 430614 513439 430616
rect 539948 430672 542419 430674
rect 539948 430616 542358 430672
rect 542414 430616 542419 430672
rect 539948 430614 542419 430616
rect 567916 430672 570019 430674
rect 567916 430616 569958 430672
rect 570014 430616 570019 430672
rect 567916 430614 570019 430616
rect 37917 430611 37983 430614
rect 66253 430611 66319 430614
rect 93853 430611 93919 430614
rect 121453 430611 121519 430614
rect 149053 430611 149119 430614
rect 178033 430611 178099 430614
rect 233233 430611 233299 430614
rect 262213 430611 262279 430614
rect 289813 430611 289879 430614
rect 317413 430611 317479 430614
rect 345013 430611 345079 430614
rect 401593 430611 401659 430614
rect 429193 430611 429259 430614
rect 458173 430611 458239 430614
rect 485773 430611 485839 430614
rect 513373 430611 513439 430614
rect 542353 430611 542419 430614
rect 569953 430611 570019 430614
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 583520 404820 584960 405060
rect 13721 404290 13787 404293
rect 42701 404290 42767 404293
rect 70301 404290 70367 404293
rect 97901 404290 97967 404293
rect 126881 404290 126947 404293
rect 154481 404290 154547 404293
rect 182081 404290 182147 404293
rect 209681 404290 209747 404293
rect 238661 404290 238727 404293
rect 266261 404290 266327 404293
rect 293861 404290 293927 404293
rect 322841 404290 322907 404293
rect 350441 404290 350507 404293
rect 378041 404290 378107 404293
rect 405641 404290 405707 404293
rect 434621 404290 434687 404293
rect 462221 404290 462287 404293
rect 489821 404290 489887 404293
rect 518801 404290 518867 404293
rect 545757 404290 545823 404293
rect 13721 404288 16100 404290
rect 13721 404232 13726 404288
rect 13782 404232 16100 404288
rect 13721 404230 16100 404232
rect 42701 404288 44068 404290
rect 42701 404232 42706 404288
rect 42762 404232 44068 404288
rect 42701 404230 44068 404232
rect 70301 404288 72036 404290
rect 70301 404232 70306 404288
rect 70362 404232 72036 404288
rect 70301 404230 72036 404232
rect 97901 404288 100188 404290
rect 97901 404232 97906 404288
rect 97962 404232 100188 404288
rect 97901 404230 100188 404232
rect 126881 404288 128156 404290
rect 126881 404232 126886 404288
rect 126942 404232 128156 404288
rect 126881 404230 128156 404232
rect 154481 404288 156124 404290
rect 154481 404232 154486 404288
rect 154542 404232 156124 404288
rect 154481 404230 156124 404232
rect 182081 404288 184092 404290
rect 182081 404232 182086 404288
rect 182142 404232 184092 404288
rect 182081 404230 184092 404232
rect 209681 404288 212060 404290
rect 209681 404232 209686 404288
rect 209742 404232 212060 404288
rect 209681 404230 212060 404232
rect 238661 404288 240212 404290
rect 238661 404232 238666 404288
rect 238722 404232 240212 404288
rect 238661 404230 240212 404232
rect 266261 404288 268180 404290
rect 266261 404232 266266 404288
rect 266322 404232 268180 404288
rect 266261 404230 268180 404232
rect 293861 404288 296148 404290
rect 293861 404232 293866 404288
rect 293922 404232 296148 404288
rect 293861 404230 296148 404232
rect 322841 404288 324116 404290
rect 322841 404232 322846 404288
rect 322902 404232 324116 404288
rect 322841 404230 324116 404232
rect 350441 404288 352084 404290
rect 350441 404232 350446 404288
rect 350502 404232 352084 404288
rect 350441 404230 352084 404232
rect 378041 404288 380052 404290
rect 378041 404232 378046 404288
rect 378102 404232 380052 404288
rect 378041 404230 380052 404232
rect 405641 404288 408204 404290
rect 405641 404232 405646 404288
rect 405702 404232 408204 404288
rect 405641 404230 408204 404232
rect 434621 404288 436172 404290
rect 434621 404232 434626 404288
rect 434682 404232 436172 404288
rect 434621 404230 436172 404232
rect 462221 404288 464140 404290
rect 462221 404232 462226 404288
rect 462282 404232 464140 404288
rect 462221 404230 464140 404232
rect 489821 404288 492108 404290
rect 489821 404232 489826 404288
rect 489882 404232 492108 404288
rect 489821 404230 492108 404232
rect 518801 404288 520076 404290
rect 518801 404232 518806 404288
rect 518862 404232 520076 404288
rect 518801 404230 520076 404232
rect 545757 404288 548044 404290
rect 545757 404232 545762 404288
rect 545818 404232 548044 404288
rect 545757 404230 548044 404232
rect 13721 404227 13787 404230
rect 42701 404227 42767 404230
rect 70301 404227 70367 404230
rect 97901 404227 97967 404230
rect 126881 404227 126947 404230
rect 154481 404227 154547 404230
rect 182081 404227 182147 404230
rect 209681 404227 209747 404230
rect 238661 404227 238727 404230
rect 266261 404227 266327 404230
rect 293861 404227 293927 404230
rect 322841 404227 322907 404230
rect 350441 404227 350507 404230
rect 378041 404227 378107 404230
rect 405641 404227 405707 404230
rect 434621 404227 434687 404230
rect 462221 404227 462287 404230
rect 489821 404227 489887 404230
rect 518801 404227 518867 404230
rect 545757 404227 545823 404230
rect 37917 403610 37983 403613
rect 66253 403610 66319 403613
rect 93853 403610 93919 403613
rect 121453 403610 121519 403613
rect 149053 403610 149119 403613
rect 178033 403610 178099 403613
rect 205633 403610 205699 403613
rect 233233 403610 233299 403613
rect 262213 403610 262279 403613
rect 289813 403610 289879 403613
rect 317413 403610 317479 403613
rect 345013 403610 345079 403613
rect 373993 403610 374059 403613
rect 401593 403610 401659 403613
rect 429193 403610 429259 403613
rect 458173 403610 458239 403613
rect 485773 403610 485839 403613
rect 513373 403610 513439 403613
rect 542353 403610 542419 403613
rect 569953 403610 570019 403613
rect 35788 403608 37983 403610
rect 35788 403552 37922 403608
rect 37978 403552 37983 403608
rect 35788 403550 37983 403552
rect 63940 403608 66319 403610
rect 63940 403552 66258 403608
rect 66314 403552 66319 403608
rect 63940 403550 66319 403552
rect 91908 403608 93919 403610
rect 91908 403552 93858 403608
rect 93914 403552 93919 403608
rect 91908 403550 93919 403552
rect 119876 403608 121519 403610
rect 119876 403552 121458 403608
rect 121514 403552 121519 403608
rect 119876 403550 121519 403552
rect 147844 403608 149119 403610
rect 147844 403552 149058 403608
rect 149114 403552 149119 403608
rect 147844 403550 149119 403552
rect 175812 403608 178099 403610
rect 175812 403552 178038 403608
rect 178094 403552 178099 403608
rect 175812 403550 178099 403552
rect 203964 403608 205699 403610
rect 203964 403552 205638 403608
rect 205694 403552 205699 403608
rect 203964 403550 205699 403552
rect 231932 403608 233299 403610
rect 231932 403552 233238 403608
rect 233294 403552 233299 403608
rect 231932 403550 233299 403552
rect 259900 403608 262279 403610
rect 259900 403552 262218 403608
rect 262274 403552 262279 403608
rect 259900 403550 262279 403552
rect 287868 403608 289879 403610
rect 287868 403552 289818 403608
rect 289874 403552 289879 403608
rect 287868 403550 289879 403552
rect 315836 403608 317479 403610
rect 315836 403552 317418 403608
rect 317474 403552 317479 403608
rect 315836 403550 317479 403552
rect 343804 403608 345079 403610
rect 343804 403552 345018 403608
rect 345074 403552 345079 403608
rect 343804 403550 345079 403552
rect 371956 403608 374059 403610
rect 371956 403552 373998 403608
rect 374054 403552 374059 403608
rect 371956 403550 374059 403552
rect 399924 403608 401659 403610
rect 399924 403552 401598 403608
rect 401654 403552 401659 403608
rect 399924 403550 401659 403552
rect 427892 403608 429259 403610
rect 427892 403552 429198 403608
rect 429254 403552 429259 403608
rect 427892 403550 429259 403552
rect 455860 403608 458239 403610
rect 455860 403552 458178 403608
rect 458234 403552 458239 403608
rect 455860 403550 458239 403552
rect 483828 403608 485839 403610
rect 483828 403552 485778 403608
rect 485834 403552 485839 403608
rect 483828 403550 485839 403552
rect 511796 403608 513439 403610
rect 511796 403552 513378 403608
rect 513434 403552 513439 403608
rect 511796 403550 513439 403552
rect 539948 403608 542419 403610
rect 539948 403552 542358 403608
rect 542414 403552 542419 403608
rect 539948 403550 542419 403552
rect 567916 403608 570019 403610
rect 567916 403552 569958 403608
rect 570014 403552 570019 403608
rect 567916 403550 570019 403552
rect 37917 403547 37983 403550
rect 66253 403547 66319 403550
rect 93853 403547 93919 403550
rect 121453 403547 121519 403550
rect 149053 403547 149119 403550
rect 178033 403547 178099 403550
rect 205633 403547 205699 403550
rect 233233 403547 233299 403550
rect 262213 403547 262279 403550
rect 289813 403547 289879 403550
rect 317413 403547 317479 403550
rect 345013 403547 345079 403550
rect 373993 403547 374059 403550
rect 401593 403547 401659 403550
rect 429193 403547 429259 403550
rect 458173 403547 458239 403550
rect 485773 403547 485839 403550
rect 513373 403547 513439 403550
rect 542353 403547 542419 403550
rect 569953 403547 570019 403550
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect 545757 377906 545823 377909
rect 545757 377904 548074 377906
rect 545757 377848 545762 377904
rect 545818 377848 548074 377904
rect 545757 377846 548074 377848
rect 545757 377843 545823 377846
rect 548014 377264 548074 377846
rect 13721 376818 13787 376821
rect 16070 376818 16130 377264
rect 13721 376816 16130 376818
rect 13721 376760 13726 376816
rect 13782 376760 16130 376816
rect 13721 376758 16130 376760
rect 42701 376818 42767 376821
rect 44038 376818 44098 377264
rect 42701 376816 44098 376818
rect 42701 376760 42706 376816
rect 42762 376760 44098 376816
rect 42701 376758 44098 376760
rect 70301 376818 70367 376821
rect 72006 376818 72066 377264
rect 70301 376816 72066 376818
rect 70301 376760 70306 376816
rect 70362 376760 72066 376816
rect 70301 376758 72066 376760
rect 97901 376818 97967 376821
rect 100158 376818 100218 377264
rect 97901 376816 100218 376818
rect 97901 376760 97906 376816
rect 97962 376760 100218 376816
rect 97901 376758 100218 376760
rect 126881 376818 126947 376821
rect 128126 376818 128186 377264
rect 126881 376816 128186 376818
rect 126881 376760 126886 376816
rect 126942 376760 128186 376816
rect 126881 376758 128186 376760
rect 154481 376818 154547 376821
rect 156094 376818 156154 377264
rect 154481 376816 156154 376818
rect 154481 376760 154486 376816
rect 154542 376760 156154 376816
rect 154481 376758 156154 376760
rect 182081 376818 182147 376821
rect 184062 376818 184122 377264
rect 209681 377090 209747 377093
rect 212030 377090 212090 377264
rect 209681 377088 212090 377090
rect 209681 377032 209686 377088
rect 209742 377032 212090 377088
rect 209681 377030 212090 377032
rect 238661 377090 238727 377093
rect 240182 377090 240242 377264
rect 238661 377088 240242 377090
rect 238661 377032 238666 377088
rect 238722 377032 240242 377088
rect 238661 377030 240242 377032
rect 266261 377090 266327 377093
rect 268150 377090 268210 377264
rect 266261 377088 268210 377090
rect 266261 377032 266266 377088
rect 266322 377032 268210 377088
rect 266261 377030 268210 377032
rect 209681 377027 209747 377030
rect 238661 377027 238727 377030
rect 266261 377027 266327 377030
rect 182081 376816 184122 376818
rect 182081 376760 182086 376816
rect 182142 376760 184122 376816
rect 182081 376758 184122 376760
rect 293861 376818 293927 376821
rect 296118 376818 296178 377264
rect 293861 376816 296178 376818
rect 293861 376760 293866 376816
rect 293922 376760 296178 376816
rect 293861 376758 296178 376760
rect 322841 376818 322907 376821
rect 324086 376818 324146 377264
rect 322841 376816 324146 376818
rect 322841 376760 322846 376816
rect 322902 376760 324146 376816
rect 322841 376758 324146 376760
rect 350441 376818 350507 376821
rect 352054 376818 352114 377264
rect 350441 376816 352114 376818
rect 350441 376760 350446 376816
rect 350502 376760 352114 376816
rect 350441 376758 352114 376760
rect 378041 376818 378107 376821
rect 380022 376818 380082 377264
rect 378041 376816 380082 376818
rect 378041 376760 378046 376816
rect 378102 376760 380082 376816
rect 378041 376758 380082 376760
rect 405641 376818 405707 376821
rect 408174 376818 408234 377264
rect 405641 376816 408234 376818
rect 405641 376760 405646 376816
rect 405702 376760 408234 376816
rect 405641 376758 408234 376760
rect 434621 376818 434687 376821
rect 436142 376818 436202 377264
rect 434621 376816 436202 376818
rect 434621 376760 434626 376816
rect 434682 376760 436202 376816
rect 434621 376758 436202 376760
rect 462221 376818 462287 376821
rect 464110 376818 464170 377264
rect 489821 377090 489887 377093
rect 492078 377090 492138 377264
rect 489821 377088 492138 377090
rect 489821 377032 489826 377088
rect 489882 377032 492138 377088
rect 489821 377030 492138 377032
rect 518801 377090 518867 377093
rect 520046 377090 520106 377264
rect 518801 377088 520106 377090
rect 518801 377032 518806 377088
rect 518862 377032 520106 377088
rect 518801 377030 520106 377032
rect 489821 377027 489887 377030
rect 518801 377027 518867 377030
rect 462221 376816 464170 376818
rect 462221 376760 462226 376816
rect 462282 376760 464170 376816
rect 462221 376758 464170 376760
rect 13721 376755 13787 376758
rect 42701 376755 42767 376758
rect 70301 376755 70367 376758
rect 97901 376755 97967 376758
rect 126881 376755 126947 376758
rect 154481 376755 154547 376758
rect 182081 376755 182147 376758
rect 293861 376755 293927 376758
rect 322841 376755 322907 376758
rect 350441 376755 350507 376758
rect 378041 376755 378107 376758
rect 405641 376755 405707 376758
rect 434621 376755 434687 376758
rect 462221 376755 462287 376758
rect 35758 376002 35818 376584
rect 37917 376002 37983 376005
rect 35758 376000 37983 376002
rect 35758 375944 37922 376000
rect 37978 375944 37983 376000
rect 35758 375942 37983 375944
rect 63910 376002 63970 376584
rect 66253 376002 66319 376005
rect 63910 376000 66319 376002
rect 63910 375944 66258 376000
rect 66314 375944 66319 376000
rect 63910 375942 66319 375944
rect 91878 376002 91938 376584
rect 93853 376002 93919 376005
rect 91878 376000 93919 376002
rect 91878 375944 93858 376000
rect 93914 375944 93919 376000
rect 91878 375942 93919 375944
rect 119846 376002 119906 376584
rect 121453 376002 121519 376005
rect 119846 376000 121519 376002
rect 119846 375944 121458 376000
rect 121514 375944 121519 376000
rect 119846 375942 121519 375944
rect 147814 376002 147874 376584
rect 149053 376002 149119 376005
rect 147814 376000 149119 376002
rect 147814 375944 149058 376000
rect 149114 375944 149119 376000
rect 147814 375942 149119 375944
rect 175782 376002 175842 376584
rect 178033 376002 178099 376005
rect 175782 376000 178099 376002
rect 175782 375944 178038 376000
rect 178094 375944 178099 376000
rect 175782 375942 178099 375944
rect 203934 376002 203994 376584
rect 205633 376002 205699 376005
rect 203934 376000 205699 376002
rect 203934 375944 205638 376000
rect 205694 375944 205699 376000
rect 203934 375942 205699 375944
rect 231902 376002 231962 376584
rect 233233 376002 233299 376005
rect 231902 376000 233299 376002
rect 231902 375944 233238 376000
rect 233294 375944 233299 376000
rect 231902 375942 233299 375944
rect 259870 376002 259930 376584
rect 260741 376002 260807 376005
rect 259870 376000 260807 376002
rect 259870 375944 260746 376000
rect 260802 375944 260807 376000
rect 259870 375942 260807 375944
rect 287838 376002 287898 376584
rect 289813 376002 289879 376005
rect 287838 376000 289879 376002
rect 287838 375944 289818 376000
rect 289874 375944 289879 376000
rect 287838 375942 289879 375944
rect 315806 376002 315866 376584
rect 317413 376002 317479 376005
rect 315806 376000 317479 376002
rect 315806 375944 317418 376000
rect 317474 375944 317479 376000
rect 315806 375942 317479 375944
rect 343774 376002 343834 376584
rect 345013 376002 345079 376005
rect 343774 376000 345079 376002
rect 343774 375944 345018 376000
rect 345074 375944 345079 376000
rect 343774 375942 345079 375944
rect 371926 376002 371986 376584
rect 373993 376002 374059 376005
rect 371926 376000 374059 376002
rect 371926 375944 373998 376000
rect 374054 375944 374059 376000
rect 371926 375942 374059 375944
rect 399894 376002 399954 376584
rect 401593 376002 401659 376005
rect 399894 376000 401659 376002
rect 399894 375944 401598 376000
rect 401654 375944 401659 376000
rect 399894 375942 401659 375944
rect 427862 376002 427922 376584
rect 429193 376002 429259 376005
rect 427862 376000 429259 376002
rect 427862 375944 429198 376000
rect 429254 375944 429259 376000
rect 427862 375942 429259 375944
rect 455830 376002 455890 376584
rect 458173 376002 458239 376005
rect 455830 376000 458239 376002
rect 455830 375944 458178 376000
rect 458234 375944 458239 376000
rect 455830 375942 458239 375944
rect 483798 376002 483858 376584
rect 485773 376002 485839 376005
rect 483798 376000 485839 376002
rect 483798 375944 485778 376000
rect 485834 375944 485839 376000
rect 483798 375942 485839 375944
rect 511766 376002 511826 376584
rect 513373 376002 513439 376005
rect 511766 376000 513439 376002
rect 511766 375944 513378 376000
rect 513434 375944 513439 376000
rect 511766 375942 513439 375944
rect 539918 376002 539978 376584
rect 540881 376002 540947 376005
rect 539918 376000 540947 376002
rect 539918 375944 540886 376000
rect 540942 375944 540947 376000
rect 539918 375942 540947 375944
rect 567886 376002 567946 376584
rect 569953 376002 570019 376005
rect 567886 376000 570019 376002
rect 567886 375944 569958 376000
rect 570014 375944 570019 376000
rect 567886 375942 570019 375944
rect 37917 375939 37983 375942
rect 66253 375939 66319 375942
rect 93853 375939 93919 375942
rect 121453 375939 121519 375942
rect 149053 375939 149119 375942
rect 178033 375939 178099 375942
rect 205633 375939 205699 375942
rect 233233 375939 233299 375942
rect 260741 375939 260807 375942
rect 289813 375939 289879 375942
rect 317413 375939 317479 375942
rect 345013 375939 345079 375942
rect 373993 375939 374059 375942
rect 401593 375939 401659 375942
rect 429193 375939 429259 375942
rect 458173 375939 458239 375942
rect 485773 375939 485839 375942
rect 513373 375939 513439 375942
rect 540881 375939 540947 375942
rect 569953 375939 570019 375942
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 583520 351780 584960 352020
rect 13721 350298 13787 350301
rect 42701 350298 42767 350301
rect 70301 350298 70367 350301
rect 97901 350298 97967 350301
rect 126881 350298 126947 350301
rect 154481 350298 154547 350301
rect 182081 350298 182147 350301
rect 209681 350298 209747 350301
rect 238661 350298 238727 350301
rect 266261 350298 266327 350301
rect 293861 350298 293927 350301
rect 322841 350298 322907 350301
rect 350441 350298 350507 350301
rect 378041 350298 378107 350301
rect 405641 350298 405707 350301
rect 434621 350298 434687 350301
rect 462221 350298 462287 350301
rect 489821 350298 489887 350301
rect 518801 350298 518867 350301
rect 545757 350298 545823 350301
rect 13721 350296 16100 350298
rect 13721 350240 13726 350296
rect 13782 350240 16100 350296
rect 13721 350238 16100 350240
rect 42701 350296 44068 350298
rect 42701 350240 42706 350296
rect 42762 350240 44068 350296
rect 42701 350238 44068 350240
rect 70301 350296 72036 350298
rect 70301 350240 70306 350296
rect 70362 350240 72036 350296
rect 70301 350238 72036 350240
rect 97901 350296 100188 350298
rect 97901 350240 97906 350296
rect 97962 350240 100188 350296
rect 97901 350238 100188 350240
rect 126881 350296 128156 350298
rect 126881 350240 126886 350296
rect 126942 350240 128156 350296
rect 126881 350238 128156 350240
rect 154481 350296 156124 350298
rect 154481 350240 154486 350296
rect 154542 350240 156124 350296
rect 154481 350238 156124 350240
rect 182081 350296 184092 350298
rect 182081 350240 182086 350296
rect 182142 350240 184092 350296
rect 182081 350238 184092 350240
rect 209681 350296 212060 350298
rect 209681 350240 209686 350296
rect 209742 350240 212060 350296
rect 209681 350238 212060 350240
rect 238661 350296 240212 350298
rect 238661 350240 238666 350296
rect 238722 350240 240212 350296
rect 238661 350238 240212 350240
rect 266261 350296 268180 350298
rect 266261 350240 266266 350296
rect 266322 350240 268180 350296
rect 266261 350238 268180 350240
rect 293861 350296 296148 350298
rect 293861 350240 293866 350296
rect 293922 350240 296148 350296
rect 293861 350238 296148 350240
rect 322841 350296 324116 350298
rect 322841 350240 322846 350296
rect 322902 350240 324116 350296
rect 322841 350238 324116 350240
rect 350441 350296 352084 350298
rect 350441 350240 350446 350296
rect 350502 350240 352084 350296
rect 350441 350238 352084 350240
rect 378041 350296 380052 350298
rect 378041 350240 378046 350296
rect 378102 350240 380052 350296
rect 378041 350238 380052 350240
rect 405641 350296 408204 350298
rect 405641 350240 405646 350296
rect 405702 350240 408204 350296
rect 405641 350238 408204 350240
rect 434621 350296 436172 350298
rect 434621 350240 434626 350296
rect 434682 350240 436172 350296
rect 434621 350238 436172 350240
rect 462221 350296 464140 350298
rect 462221 350240 462226 350296
rect 462282 350240 464140 350296
rect 462221 350238 464140 350240
rect 489821 350296 492108 350298
rect 489821 350240 489826 350296
rect 489882 350240 492108 350296
rect 489821 350238 492108 350240
rect 518801 350296 520076 350298
rect 518801 350240 518806 350296
rect 518862 350240 520076 350296
rect 518801 350238 520076 350240
rect 545757 350296 548044 350298
rect 545757 350240 545762 350296
rect 545818 350240 548044 350296
rect 545757 350238 548044 350240
rect 13721 350235 13787 350238
rect 42701 350235 42767 350238
rect 70301 350235 70367 350238
rect 97901 350235 97967 350238
rect 126881 350235 126947 350238
rect 154481 350235 154547 350238
rect 182081 350235 182147 350238
rect 209681 350235 209747 350238
rect 238661 350235 238727 350238
rect 266261 350235 266327 350238
rect 293861 350235 293927 350238
rect 322841 350235 322907 350238
rect 350441 350235 350507 350238
rect 378041 350235 378107 350238
rect 405641 350235 405707 350238
rect 434621 350235 434687 350238
rect 462221 350235 462287 350238
rect 489821 350235 489887 350238
rect 518801 350235 518867 350238
rect 545757 350235 545823 350238
rect 37917 349618 37983 349621
rect 66253 349618 66319 349621
rect 93853 349618 93919 349621
rect 121453 349618 121519 349621
rect 149053 349618 149119 349621
rect 178033 349618 178099 349621
rect 205633 349618 205699 349621
rect 233233 349618 233299 349621
rect 262213 349618 262279 349621
rect 289813 349618 289879 349621
rect 317413 349618 317479 349621
rect 345013 349618 345079 349621
rect 373993 349618 374059 349621
rect 401593 349618 401659 349621
rect 429193 349618 429259 349621
rect 458173 349618 458239 349621
rect 485773 349618 485839 349621
rect 513373 349618 513439 349621
rect 542353 349618 542419 349621
rect 569953 349618 570019 349621
rect 35788 349616 37983 349618
rect 35788 349560 37922 349616
rect 37978 349560 37983 349616
rect 35788 349558 37983 349560
rect 63940 349616 66319 349618
rect 63940 349560 66258 349616
rect 66314 349560 66319 349616
rect 63940 349558 66319 349560
rect 91908 349616 93919 349618
rect 91908 349560 93858 349616
rect 93914 349560 93919 349616
rect 91908 349558 93919 349560
rect 119876 349616 121519 349618
rect 119876 349560 121458 349616
rect 121514 349560 121519 349616
rect 119876 349558 121519 349560
rect 147844 349616 149119 349618
rect 147844 349560 149058 349616
rect 149114 349560 149119 349616
rect 147844 349558 149119 349560
rect 175812 349616 178099 349618
rect 175812 349560 178038 349616
rect 178094 349560 178099 349616
rect 175812 349558 178099 349560
rect 203964 349616 205699 349618
rect 203964 349560 205638 349616
rect 205694 349560 205699 349616
rect 203964 349558 205699 349560
rect 231932 349616 233299 349618
rect 231932 349560 233238 349616
rect 233294 349560 233299 349616
rect 231932 349558 233299 349560
rect 259900 349616 262279 349618
rect 259900 349560 262218 349616
rect 262274 349560 262279 349616
rect 259900 349558 262279 349560
rect 287868 349616 289879 349618
rect 287868 349560 289818 349616
rect 289874 349560 289879 349616
rect 287868 349558 289879 349560
rect 315836 349616 317479 349618
rect 315836 349560 317418 349616
rect 317474 349560 317479 349616
rect 315836 349558 317479 349560
rect 343804 349616 345079 349618
rect 343804 349560 345018 349616
rect 345074 349560 345079 349616
rect 343804 349558 345079 349560
rect 371956 349616 374059 349618
rect 371956 349560 373998 349616
rect 374054 349560 374059 349616
rect 371956 349558 374059 349560
rect 399924 349616 401659 349618
rect 399924 349560 401598 349616
rect 401654 349560 401659 349616
rect 399924 349558 401659 349560
rect 427892 349616 429259 349618
rect 427892 349560 429198 349616
rect 429254 349560 429259 349616
rect 427892 349558 429259 349560
rect 455860 349616 458239 349618
rect 455860 349560 458178 349616
rect 458234 349560 458239 349616
rect 455860 349558 458239 349560
rect 483828 349616 485839 349618
rect 483828 349560 485778 349616
rect 485834 349560 485839 349616
rect 483828 349558 485839 349560
rect 511796 349616 513439 349618
rect 511796 349560 513378 349616
rect 513434 349560 513439 349616
rect 511796 349558 513439 349560
rect 539948 349616 542419 349618
rect 539948 349560 542358 349616
rect 542414 349560 542419 349616
rect 539948 349558 542419 349560
rect 567916 349616 570019 349618
rect 567916 349560 569958 349616
rect 570014 349560 570019 349616
rect 567916 349558 570019 349560
rect 37917 349555 37983 349558
rect 66253 349555 66319 349558
rect 93853 349555 93919 349558
rect 121453 349555 121519 349558
rect 149053 349555 149119 349558
rect 178033 349555 178099 349558
rect 205633 349555 205699 349558
rect 233233 349555 233299 349558
rect 262213 349555 262279 349558
rect 289813 349555 289879 349558
rect 317413 349555 317479 349558
rect 345013 349555 345079 349558
rect 373993 349555 374059 349558
rect 401593 349555 401659 349558
rect 429193 349555 429259 349558
rect 458173 349555 458239 349558
rect 485773 349555 485839 349558
rect 513373 349555 513439 349558
rect 542353 349555 542419 349558
rect 569953 349555 570019 349558
rect -960 345402 480 345492
rect 3601 345402 3667 345405
rect -960 345400 3667 345402
rect -960 345344 3606 345400
rect 3662 345344 3667 345400
rect -960 345342 3667 345344
rect -960 345252 480 345342
rect 3601 345339 3667 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect 209681 323914 209747 323917
rect 266261 323914 266327 323917
rect 405641 323914 405707 323917
rect 462221 323914 462287 323917
rect 545757 323914 545823 323917
rect 209681 323912 212090 323914
rect 209681 323856 209686 323912
rect 209742 323856 212090 323912
rect 209681 323854 212090 323856
rect 209681 323851 209747 323854
rect 212030 323272 212090 323854
rect 266261 323912 268210 323914
rect 266261 323856 266266 323912
rect 266322 323856 268210 323912
rect 266261 323854 268210 323856
rect 266261 323851 266327 323854
rect 268150 323272 268210 323854
rect 405641 323912 408234 323914
rect 405641 323856 405646 323912
rect 405702 323856 408234 323912
rect 405641 323854 408234 323856
rect 405641 323851 405707 323854
rect 408174 323272 408234 323854
rect 462221 323912 464170 323914
rect 462221 323856 462226 323912
rect 462282 323856 464170 323912
rect 462221 323854 464170 323856
rect 462221 323851 462287 323854
rect 464110 323272 464170 323854
rect 545757 323912 548074 323914
rect 545757 323856 545762 323912
rect 545818 323856 548074 323912
rect 545757 323854 548074 323856
rect 545757 323851 545823 323854
rect 548014 323272 548074 323854
rect 13721 322962 13787 322965
rect 16070 322962 16130 323272
rect 13721 322960 16130 322962
rect 13721 322904 13726 322960
rect 13782 322904 16130 322960
rect 13721 322902 16130 322904
rect 42701 322962 42767 322965
rect 44038 322962 44098 323272
rect 42701 322960 44098 322962
rect 42701 322904 42706 322960
rect 42762 322904 44098 322960
rect 42701 322902 44098 322904
rect 70301 322962 70367 322965
rect 72006 322962 72066 323272
rect 70301 322960 72066 322962
rect 70301 322904 70306 322960
rect 70362 322904 72066 322960
rect 70301 322902 72066 322904
rect 97901 322962 97967 322965
rect 100158 322962 100218 323272
rect 97901 322960 100218 322962
rect 97901 322904 97906 322960
rect 97962 322904 100218 322960
rect 97901 322902 100218 322904
rect 126881 322962 126947 322965
rect 128126 322962 128186 323272
rect 126881 322960 128186 322962
rect 126881 322904 126886 322960
rect 126942 322904 128186 322960
rect 126881 322902 128186 322904
rect 154481 322962 154547 322965
rect 156094 322962 156154 323272
rect 154481 322960 156154 322962
rect 154481 322904 154486 322960
rect 154542 322904 156154 322960
rect 154481 322902 156154 322904
rect 182081 322962 182147 322965
rect 184062 322962 184122 323272
rect 182081 322960 184122 322962
rect 182081 322904 182086 322960
rect 182142 322904 184122 322960
rect 182081 322902 184122 322904
rect 238661 322962 238727 322965
rect 240182 322962 240242 323272
rect 238661 322960 240242 322962
rect 238661 322904 238666 322960
rect 238722 322904 240242 322960
rect 238661 322902 240242 322904
rect 293861 322962 293927 322965
rect 296118 322962 296178 323272
rect 293861 322960 296178 322962
rect 293861 322904 293866 322960
rect 293922 322904 296178 322960
rect 293861 322902 296178 322904
rect 322841 322962 322907 322965
rect 324086 322962 324146 323272
rect 322841 322960 324146 322962
rect 322841 322904 322846 322960
rect 322902 322904 324146 322960
rect 322841 322902 324146 322904
rect 350441 322962 350507 322965
rect 352054 322962 352114 323272
rect 350441 322960 352114 322962
rect 350441 322904 350446 322960
rect 350502 322904 352114 322960
rect 350441 322902 352114 322904
rect 378041 322962 378107 322965
rect 380022 322962 380082 323272
rect 378041 322960 380082 322962
rect 378041 322904 378046 322960
rect 378102 322904 380082 322960
rect 378041 322902 380082 322904
rect 434621 322962 434687 322965
rect 436142 322962 436202 323272
rect 434621 322960 436202 322962
rect 434621 322904 434626 322960
rect 434682 322904 436202 322960
rect 434621 322902 436202 322904
rect 489821 322962 489887 322965
rect 492078 322962 492138 323272
rect 489821 322960 492138 322962
rect 489821 322904 489826 322960
rect 489882 322904 492138 322960
rect 489821 322902 492138 322904
rect 518801 322962 518867 322965
rect 520046 322962 520106 323272
rect 518801 322960 520106 322962
rect 518801 322904 518806 322960
rect 518862 322904 520106 322960
rect 518801 322902 520106 322904
rect 13721 322899 13787 322902
rect 42701 322899 42767 322902
rect 70301 322899 70367 322902
rect 97901 322899 97967 322902
rect 126881 322899 126947 322902
rect 154481 322899 154547 322902
rect 182081 322899 182147 322902
rect 238661 322899 238727 322902
rect 293861 322899 293927 322902
rect 322841 322899 322907 322902
rect 350441 322899 350507 322902
rect 378041 322899 378107 322902
rect 434621 322899 434687 322902
rect 489821 322899 489887 322902
rect 518801 322899 518867 322902
rect 262213 322826 262279 322829
rect 317413 322826 317479 322829
rect 458173 322826 458239 322829
rect 513373 322826 513439 322829
rect 259870 322824 262279 322826
rect 259870 322768 262218 322824
rect 262274 322768 262279 322824
rect 259870 322766 262279 322768
rect 259870 322592 259930 322766
rect 262213 322763 262279 322766
rect 315806 322824 317479 322826
rect 315806 322768 317418 322824
rect 317474 322768 317479 322824
rect 315806 322766 317479 322768
rect 315806 322592 315866 322766
rect 317413 322763 317479 322766
rect 455830 322824 458239 322826
rect 455830 322768 458178 322824
rect 458234 322768 458239 322824
rect 455830 322766 458239 322768
rect 455830 322592 455890 322766
rect 458173 322763 458239 322766
rect 511766 322824 513439 322826
rect 511766 322768 513378 322824
rect 513434 322768 513439 322824
rect 511766 322766 513439 322768
rect 511766 322592 511826 322766
rect 513373 322763 513439 322766
rect 35758 322010 35818 322592
rect 37917 322010 37983 322013
rect 35758 322008 37983 322010
rect 35758 321952 37922 322008
rect 37978 321952 37983 322008
rect 35758 321950 37983 321952
rect 63910 322010 63970 322592
rect 66253 322010 66319 322013
rect 63910 322008 66319 322010
rect 63910 321952 66258 322008
rect 66314 321952 66319 322008
rect 63910 321950 66319 321952
rect 91878 322010 91938 322592
rect 93853 322010 93919 322013
rect 91878 322008 93919 322010
rect 91878 321952 93858 322008
rect 93914 321952 93919 322008
rect 91878 321950 93919 321952
rect 119846 322010 119906 322592
rect 121453 322010 121519 322013
rect 119846 322008 121519 322010
rect 119846 321952 121458 322008
rect 121514 321952 121519 322008
rect 119846 321950 121519 321952
rect 147814 322010 147874 322592
rect 149053 322010 149119 322013
rect 147814 322008 149119 322010
rect 147814 321952 149058 322008
rect 149114 321952 149119 322008
rect 147814 321950 149119 321952
rect 175782 322010 175842 322592
rect 178033 322010 178099 322013
rect 175782 322008 178099 322010
rect 175782 321952 178038 322008
rect 178094 321952 178099 322008
rect 175782 321950 178099 321952
rect 203934 322010 203994 322592
rect 205633 322010 205699 322013
rect 203934 322008 205699 322010
rect 203934 321952 205638 322008
rect 205694 321952 205699 322008
rect 203934 321950 205699 321952
rect 231902 322010 231962 322592
rect 233233 322010 233299 322013
rect 231902 322008 233299 322010
rect 231902 321952 233238 322008
rect 233294 321952 233299 322008
rect 231902 321950 233299 321952
rect 287838 322010 287898 322592
rect 289813 322010 289879 322013
rect 287838 322008 289879 322010
rect 287838 321952 289818 322008
rect 289874 321952 289879 322008
rect 287838 321950 289879 321952
rect 343774 322010 343834 322592
rect 345013 322010 345079 322013
rect 343774 322008 345079 322010
rect 343774 321952 345018 322008
rect 345074 321952 345079 322008
rect 343774 321950 345079 321952
rect 371926 322010 371986 322592
rect 373993 322010 374059 322013
rect 371926 322008 374059 322010
rect 371926 321952 373998 322008
rect 374054 321952 374059 322008
rect 371926 321950 374059 321952
rect 399894 322010 399954 322592
rect 401593 322010 401659 322013
rect 399894 322008 401659 322010
rect 399894 321952 401598 322008
rect 401654 321952 401659 322008
rect 399894 321950 401659 321952
rect 427862 322010 427922 322592
rect 429193 322010 429259 322013
rect 427862 322008 429259 322010
rect 427862 321952 429198 322008
rect 429254 321952 429259 322008
rect 427862 321950 429259 321952
rect 483798 322010 483858 322592
rect 485773 322010 485839 322013
rect 483798 322008 485839 322010
rect 483798 321952 485778 322008
rect 485834 321952 485839 322008
rect 483798 321950 485839 321952
rect 539918 322010 539978 322592
rect 542353 322010 542419 322013
rect 539918 322008 542419 322010
rect 539918 321952 542358 322008
rect 542414 321952 542419 322008
rect 539918 321950 542419 321952
rect 567886 322010 567946 322592
rect 569953 322010 570019 322013
rect 567886 322008 570019 322010
rect 567886 321952 569958 322008
rect 570014 321952 570019 322008
rect 567886 321950 570019 321952
rect 37917 321947 37983 321950
rect 66253 321947 66319 321950
rect 93853 321947 93919 321950
rect 121453 321947 121519 321950
rect 149053 321947 149119 321950
rect 178033 321947 178099 321950
rect 205633 321947 205699 321950
rect 233233 321947 233299 321950
rect 289813 321947 289879 321950
rect 345013 321947 345079 321950
rect 373993 321947 374059 321950
rect 401593 321947 401659 321950
rect 429193 321947 429259 321950
rect 485773 321947 485839 321950
rect 542353 321947 542419 321950
rect 569953 321947 570019 321950
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306234 480 306324
rect 3049 306234 3115 306237
rect -960 306232 3115 306234
rect -960 306176 3054 306232
rect 3110 306176 3115 306232
rect -960 306174 3115 306176
rect -960 306084 480 306174
rect 3049 306171 3115 306174
rect 583520 298604 584960 298844
rect 13721 296306 13787 296309
rect 42701 296306 42767 296309
rect 70301 296306 70367 296309
rect 97901 296306 97967 296309
rect 126881 296306 126947 296309
rect 154481 296306 154547 296309
rect 182081 296306 182147 296309
rect 209681 296306 209747 296309
rect 238661 296306 238727 296309
rect 266261 296306 266327 296309
rect 293861 296306 293927 296309
rect 322841 296306 322907 296309
rect 350441 296306 350507 296309
rect 378041 296306 378107 296309
rect 405641 296306 405707 296309
rect 434621 296306 434687 296309
rect 462221 296306 462287 296309
rect 489821 296306 489887 296309
rect 518801 296306 518867 296309
rect 545757 296306 545823 296309
rect 13721 296304 16100 296306
rect 13721 296248 13726 296304
rect 13782 296248 16100 296304
rect 13721 296246 16100 296248
rect 42701 296304 44068 296306
rect 42701 296248 42706 296304
rect 42762 296248 44068 296304
rect 42701 296246 44068 296248
rect 70301 296304 72036 296306
rect 70301 296248 70306 296304
rect 70362 296248 72036 296304
rect 70301 296246 72036 296248
rect 97901 296304 100188 296306
rect 97901 296248 97906 296304
rect 97962 296248 100188 296304
rect 97901 296246 100188 296248
rect 126881 296304 128156 296306
rect 126881 296248 126886 296304
rect 126942 296248 128156 296304
rect 126881 296246 128156 296248
rect 154481 296304 156124 296306
rect 154481 296248 154486 296304
rect 154542 296248 156124 296304
rect 154481 296246 156124 296248
rect 182081 296304 184092 296306
rect 182081 296248 182086 296304
rect 182142 296248 184092 296304
rect 182081 296246 184092 296248
rect 209681 296304 212060 296306
rect 209681 296248 209686 296304
rect 209742 296248 212060 296304
rect 209681 296246 212060 296248
rect 238661 296304 240212 296306
rect 238661 296248 238666 296304
rect 238722 296248 240212 296304
rect 238661 296246 240212 296248
rect 266261 296304 268180 296306
rect 266261 296248 266266 296304
rect 266322 296248 268180 296304
rect 266261 296246 268180 296248
rect 293861 296304 296148 296306
rect 293861 296248 293866 296304
rect 293922 296248 296148 296304
rect 293861 296246 296148 296248
rect 322841 296304 324116 296306
rect 322841 296248 322846 296304
rect 322902 296248 324116 296304
rect 322841 296246 324116 296248
rect 350441 296304 352084 296306
rect 350441 296248 350446 296304
rect 350502 296248 352084 296304
rect 350441 296246 352084 296248
rect 378041 296304 380052 296306
rect 378041 296248 378046 296304
rect 378102 296248 380052 296304
rect 378041 296246 380052 296248
rect 405641 296304 408204 296306
rect 405641 296248 405646 296304
rect 405702 296248 408204 296304
rect 405641 296246 408204 296248
rect 434621 296304 436172 296306
rect 434621 296248 434626 296304
rect 434682 296248 436172 296304
rect 434621 296246 436172 296248
rect 462221 296304 464140 296306
rect 462221 296248 462226 296304
rect 462282 296248 464140 296304
rect 462221 296246 464140 296248
rect 489821 296304 492108 296306
rect 489821 296248 489826 296304
rect 489882 296248 492108 296304
rect 489821 296246 492108 296248
rect 518801 296304 520076 296306
rect 518801 296248 518806 296304
rect 518862 296248 520076 296304
rect 518801 296246 520076 296248
rect 545757 296304 548044 296306
rect 545757 296248 545762 296304
rect 545818 296248 548044 296304
rect 545757 296246 548044 296248
rect 13721 296243 13787 296246
rect 42701 296243 42767 296246
rect 70301 296243 70367 296246
rect 97901 296243 97967 296246
rect 126881 296243 126947 296246
rect 154481 296243 154547 296246
rect 182081 296243 182147 296246
rect 209681 296243 209747 296246
rect 238661 296243 238727 296246
rect 266261 296243 266327 296246
rect 293861 296243 293927 296246
rect 322841 296243 322907 296246
rect 350441 296243 350507 296246
rect 378041 296243 378107 296246
rect 405641 296243 405707 296246
rect 434621 296243 434687 296246
rect 462221 296243 462287 296246
rect 489821 296243 489887 296246
rect 518801 296243 518867 296246
rect 545757 296243 545823 296246
rect 37917 295626 37983 295629
rect 66253 295626 66319 295629
rect 93853 295626 93919 295629
rect 121453 295626 121519 295629
rect 149053 295626 149119 295629
rect 178033 295626 178099 295629
rect 205633 295626 205699 295629
rect 233233 295626 233299 295629
rect 262213 295626 262279 295629
rect 289813 295626 289879 295629
rect 317413 295626 317479 295629
rect 345013 295626 345079 295629
rect 373993 295626 374059 295629
rect 401593 295626 401659 295629
rect 429193 295626 429259 295629
rect 458173 295626 458239 295629
rect 485773 295626 485839 295629
rect 513373 295626 513439 295629
rect 542353 295626 542419 295629
rect 569953 295626 570019 295629
rect 35788 295624 37983 295626
rect 35788 295568 37922 295624
rect 37978 295568 37983 295624
rect 35788 295566 37983 295568
rect 63940 295624 66319 295626
rect 63940 295568 66258 295624
rect 66314 295568 66319 295624
rect 63940 295566 66319 295568
rect 91908 295624 93919 295626
rect 91908 295568 93858 295624
rect 93914 295568 93919 295624
rect 91908 295566 93919 295568
rect 119876 295624 121519 295626
rect 119876 295568 121458 295624
rect 121514 295568 121519 295624
rect 119876 295566 121519 295568
rect 147844 295624 149119 295626
rect 147844 295568 149058 295624
rect 149114 295568 149119 295624
rect 147844 295566 149119 295568
rect 175812 295624 178099 295626
rect 175812 295568 178038 295624
rect 178094 295568 178099 295624
rect 175812 295566 178099 295568
rect 203964 295624 205699 295626
rect 203964 295568 205638 295624
rect 205694 295568 205699 295624
rect 203964 295566 205699 295568
rect 231932 295624 233299 295626
rect 231932 295568 233238 295624
rect 233294 295568 233299 295624
rect 231932 295566 233299 295568
rect 259900 295624 262279 295626
rect 259900 295568 262218 295624
rect 262274 295568 262279 295624
rect 259900 295566 262279 295568
rect 287868 295624 289879 295626
rect 287868 295568 289818 295624
rect 289874 295568 289879 295624
rect 287868 295566 289879 295568
rect 315836 295624 317479 295626
rect 315836 295568 317418 295624
rect 317474 295568 317479 295624
rect 315836 295566 317479 295568
rect 343804 295624 345079 295626
rect 343804 295568 345018 295624
rect 345074 295568 345079 295624
rect 343804 295566 345079 295568
rect 371956 295624 374059 295626
rect 371956 295568 373998 295624
rect 374054 295568 374059 295624
rect 371956 295566 374059 295568
rect 399924 295624 401659 295626
rect 399924 295568 401598 295624
rect 401654 295568 401659 295624
rect 399924 295566 401659 295568
rect 427892 295624 429259 295626
rect 427892 295568 429198 295624
rect 429254 295568 429259 295624
rect 427892 295566 429259 295568
rect 455860 295624 458239 295626
rect 455860 295568 458178 295624
rect 458234 295568 458239 295624
rect 455860 295566 458239 295568
rect 483828 295624 485839 295626
rect 483828 295568 485778 295624
rect 485834 295568 485839 295624
rect 483828 295566 485839 295568
rect 511796 295624 513439 295626
rect 511796 295568 513378 295624
rect 513434 295568 513439 295624
rect 511796 295566 513439 295568
rect 539948 295624 542419 295626
rect 539948 295568 542358 295624
rect 542414 295568 542419 295624
rect 539948 295566 542419 295568
rect 567916 295624 570019 295626
rect 567916 295568 569958 295624
rect 570014 295568 570019 295624
rect 567916 295566 570019 295568
rect 37917 295563 37983 295566
rect 66253 295563 66319 295566
rect 93853 295563 93919 295566
rect 121453 295563 121519 295566
rect 149053 295563 149119 295566
rect 178033 295563 178099 295566
rect 205633 295563 205699 295566
rect 233233 295563 233299 295566
rect 262213 295563 262279 295566
rect 289813 295563 289879 295566
rect 317413 295563 317479 295566
rect 345013 295563 345079 295566
rect 373993 295563 374059 295566
rect 401593 295563 401659 295566
rect 429193 295563 429259 295566
rect 458173 295563 458239 295566
rect 485773 295563 485839 295566
rect 513373 295563 513439 295566
rect 542353 295563 542419 295566
rect 569953 295563 570019 295566
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect 70301 269786 70367 269789
rect 545757 269786 545823 269789
rect 70301 269784 72066 269786
rect 70301 269728 70306 269784
rect 70362 269728 72066 269784
rect 70301 269726 72066 269728
rect 70301 269723 70367 269726
rect 13721 269242 13787 269245
rect 42701 269242 42767 269245
rect 13721 269240 16100 269242
rect 13721 269184 13726 269240
rect 13782 269184 16100 269240
rect 13721 269182 16100 269184
rect 42701 269240 44068 269242
rect 42701 269184 42706 269240
rect 42762 269184 44068 269240
rect 72006 269212 72066 269726
rect 545757 269784 548074 269786
rect 545757 269728 545762 269784
rect 545818 269728 548074 269784
rect 545757 269726 548074 269728
rect 545757 269723 545823 269726
rect 97901 269242 97967 269245
rect 126881 269242 126947 269245
rect 154481 269242 154547 269245
rect 182081 269242 182147 269245
rect 209681 269242 209747 269245
rect 238661 269242 238727 269245
rect 266261 269242 266327 269245
rect 293861 269242 293927 269245
rect 322841 269242 322907 269245
rect 350441 269242 350507 269245
rect 378041 269242 378107 269245
rect 405641 269242 405707 269245
rect 434621 269242 434687 269245
rect 462221 269242 462287 269245
rect 489821 269242 489887 269245
rect 518801 269242 518867 269245
rect 97901 269240 100188 269242
rect 42701 269182 44068 269184
rect 97901 269184 97906 269240
rect 97962 269184 100188 269240
rect 97901 269182 100188 269184
rect 126881 269240 128156 269242
rect 126881 269184 126886 269240
rect 126942 269184 128156 269240
rect 126881 269182 128156 269184
rect 154481 269240 156124 269242
rect 154481 269184 154486 269240
rect 154542 269184 156124 269240
rect 154481 269182 156124 269184
rect 182081 269240 184092 269242
rect 182081 269184 182086 269240
rect 182142 269184 184092 269240
rect 182081 269182 184092 269184
rect 209681 269240 212060 269242
rect 209681 269184 209686 269240
rect 209742 269184 212060 269240
rect 209681 269182 212060 269184
rect 238661 269240 240212 269242
rect 238661 269184 238666 269240
rect 238722 269184 240212 269240
rect 238661 269182 240212 269184
rect 266261 269240 268180 269242
rect 266261 269184 266266 269240
rect 266322 269184 268180 269240
rect 266261 269182 268180 269184
rect 293861 269240 296148 269242
rect 293861 269184 293866 269240
rect 293922 269184 296148 269240
rect 293861 269182 296148 269184
rect 322841 269240 324116 269242
rect 322841 269184 322846 269240
rect 322902 269184 324116 269240
rect 322841 269182 324116 269184
rect 350441 269240 352084 269242
rect 350441 269184 350446 269240
rect 350502 269184 352084 269240
rect 350441 269182 352084 269184
rect 378041 269240 380052 269242
rect 378041 269184 378046 269240
rect 378102 269184 380052 269240
rect 378041 269182 380052 269184
rect 405641 269240 408204 269242
rect 405641 269184 405646 269240
rect 405702 269184 408204 269240
rect 405641 269182 408204 269184
rect 434621 269240 436172 269242
rect 434621 269184 434626 269240
rect 434682 269184 436172 269240
rect 434621 269182 436172 269184
rect 462221 269240 464140 269242
rect 462221 269184 462226 269240
rect 462282 269184 464140 269240
rect 462221 269182 464140 269184
rect 489821 269240 492108 269242
rect 489821 269184 489826 269240
rect 489882 269184 492108 269240
rect 489821 269182 492108 269184
rect 518801 269240 520076 269242
rect 518801 269184 518806 269240
rect 518862 269184 520076 269240
rect 548014 269212 548074 269726
rect 518801 269182 520076 269184
rect 13721 269179 13787 269182
rect 42701 269179 42767 269182
rect 97901 269179 97967 269182
rect 126881 269179 126947 269182
rect 154481 269179 154547 269182
rect 182081 269179 182147 269182
rect 209681 269179 209747 269182
rect 238661 269179 238727 269182
rect 266261 269179 266327 269182
rect 293861 269179 293927 269182
rect 322841 269179 322907 269182
rect 350441 269179 350507 269182
rect 378041 269179 378107 269182
rect 405641 269179 405707 269182
rect 434621 269179 434687 269182
rect 462221 269179 462287 269182
rect 489821 269179 489887 269182
rect 518801 269179 518867 269182
rect 205633 269106 205699 269109
rect 373993 269106 374059 269109
rect 203934 269104 205699 269106
rect 203934 269048 205638 269104
rect 205694 269048 205699 269104
rect 203934 269046 205699 269048
rect 37917 268562 37983 268565
rect 66253 268562 66319 268565
rect 93853 268562 93919 268565
rect 121453 268562 121519 268565
rect 149053 268562 149119 268565
rect 178033 268562 178099 268565
rect 35788 268560 37983 268562
rect 35788 268504 37922 268560
rect 37978 268504 37983 268560
rect 35788 268502 37983 268504
rect 63940 268560 66319 268562
rect 63940 268504 66258 268560
rect 66314 268504 66319 268560
rect 63940 268502 66319 268504
rect 91908 268560 93919 268562
rect 91908 268504 93858 268560
rect 93914 268504 93919 268560
rect 91908 268502 93919 268504
rect 119876 268560 121519 268562
rect 119876 268504 121458 268560
rect 121514 268504 121519 268560
rect 119876 268502 121519 268504
rect 147844 268560 149119 268562
rect 147844 268504 149058 268560
rect 149114 268504 149119 268560
rect 147844 268502 149119 268504
rect 175812 268560 178099 268562
rect 175812 268504 178038 268560
rect 178094 268504 178099 268560
rect 203934 268532 203994 269046
rect 205633 269043 205699 269046
rect 371926 269104 374059 269106
rect 371926 269048 373998 269104
rect 374054 269048 374059 269104
rect 371926 269046 374059 269048
rect 233233 268562 233299 268565
rect 262213 268562 262279 268565
rect 289813 268562 289879 268565
rect 317413 268562 317479 268565
rect 345013 268562 345079 268565
rect 231932 268560 233299 268562
rect 175812 268502 178099 268504
rect 231932 268504 233238 268560
rect 233294 268504 233299 268560
rect 231932 268502 233299 268504
rect 259900 268560 262279 268562
rect 259900 268504 262218 268560
rect 262274 268504 262279 268560
rect 259900 268502 262279 268504
rect 287868 268560 289879 268562
rect 287868 268504 289818 268560
rect 289874 268504 289879 268560
rect 287868 268502 289879 268504
rect 315836 268560 317479 268562
rect 315836 268504 317418 268560
rect 317474 268504 317479 268560
rect 315836 268502 317479 268504
rect 343804 268560 345079 268562
rect 343804 268504 345018 268560
rect 345074 268504 345079 268560
rect 371926 268532 371986 269046
rect 373993 269043 374059 269046
rect 401593 268562 401659 268565
rect 429193 268562 429259 268565
rect 458173 268562 458239 268565
rect 485773 268562 485839 268565
rect 513373 268562 513439 268565
rect 542353 268562 542419 268565
rect 569953 268562 570019 268565
rect 399924 268560 401659 268562
rect 343804 268502 345079 268504
rect 399924 268504 401598 268560
rect 401654 268504 401659 268560
rect 399924 268502 401659 268504
rect 427892 268560 429259 268562
rect 427892 268504 429198 268560
rect 429254 268504 429259 268560
rect 427892 268502 429259 268504
rect 455860 268560 458239 268562
rect 455860 268504 458178 268560
rect 458234 268504 458239 268560
rect 455860 268502 458239 268504
rect 483828 268560 485839 268562
rect 483828 268504 485778 268560
rect 485834 268504 485839 268560
rect 483828 268502 485839 268504
rect 511796 268560 513439 268562
rect 511796 268504 513378 268560
rect 513434 268504 513439 268560
rect 511796 268502 513439 268504
rect 539948 268560 542419 268562
rect 539948 268504 542358 268560
rect 542414 268504 542419 268560
rect 539948 268502 542419 268504
rect 567916 268560 570019 268562
rect 567916 268504 569958 268560
rect 570014 268504 570019 268560
rect 567916 268502 570019 268504
rect 37917 268499 37983 268502
rect 66253 268499 66319 268502
rect 93853 268499 93919 268502
rect 121453 268499 121519 268502
rect 149053 268499 149119 268502
rect 178033 268499 178099 268502
rect 233233 268499 233299 268502
rect 262213 268499 262279 268502
rect 289813 268499 289879 268502
rect 317413 268499 317479 268502
rect 345013 268499 345079 268502
rect 401593 268499 401659 268502
rect 429193 268499 429259 268502
rect 458173 268499 458239 268502
rect 485773 268499 485839 268502
rect 513373 268499 513439 268502
rect 542353 268499 542419 268502
rect 569953 268499 570019 268502
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 583520 245428 584960 245668
rect 13721 242314 13787 242317
rect 42701 242314 42767 242317
rect 70301 242314 70367 242317
rect 97901 242314 97967 242317
rect 126881 242314 126947 242317
rect 154481 242314 154547 242317
rect 182081 242314 182147 242317
rect 209681 242314 209747 242317
rect 238661 242314 238727 242317
rect 266261 242314 266327 242317
rect 293861 242314 293927 242317
rect 322841 242314 322907 242317
rect 350441 242314 350507 242317
rect 378041 242314 378107 242317
rect 405641 242314 405707 242317
rect 434621 242314 434687 242317
rect 462221 242314 462287 242317
rect 489821 242314 489887 242317
rect 518801 242314 518867 242317
rect 545757 242314 545823 242317
rect 13721 242312 16100 242314
rect 13721 242256 13726 242312
rect 13782 242256 16100 242312
rect 13721 242254 16100 242256
rect 42701 242312 44068 242314
rect 42701 242256 42706 242312
rect 42762 242256 44068 242312
rect 42701 242254 44068 242256
rect 70301 242312 72036 242314
rect 70301 242256 70306 242312
rect 70362 242256 72036 242312
rect 70301 242254 72036 242256
rect 97901 242312 100188 242314
rect 97901 242256 97906 242312
rect 97962 242256 100188 242312
rect 97901 242254 100188 242256
rect 126881 242312 128156 242314
rect 126881 242256 126886 242312
rect 126942 242256 128156 242312
rect 126881 242254 128156 242256
rect 154481 242312 156124 242314
rect 154481 242256 154486 242312
rect 154542 242256 156124 242312
rect 154481 242254 156124 242256
rect 182081 242312 184092 242314
rect 182081 242256 182086 242312
rect 182142 242256 184092 242312
rect 182081 242254 184092 242256
rect 209681 242312 212060 242314
rect 209681 242256 209686 242312
rect 209742 242256 212060 242312
rect 209681 242254 212060 242256
rect 238661 242312 240212 242314
rect 238661 242256 238666 242312
rect 238722 242256 240212 242312
rect 238661 242254 240212 242256
rect 266261 242312 268180 242314
rect 266261 242256 266266 242312
rect 266322 242256 268180 242312
rect 266261 242254 268180 242256
rect 293861 242312 296148 242314
rect 293861 242256 293866 242312
rect 293922 242256 296148 242312
rect 293861 242254 296148 242256
rect 322841 242312 324116 242314
rect 322841 242256 322846 242312
rect 322902 242256 324116 242312
rect 322841 242254 324116 242256
rect 350441 242312 352084 242314
rect 350441 242256 350446 242312
rect 350502 242256 352084 242312
rect 350441 242254 352084 242256
rect 378041 242312 380052 242314
rect 378041 242256 378046 242312
rect 378102 242256 380052 242312
rect 378041 242254 380052 242256
rect 405641 242312 408204 242314
rect 405641 242256 405646 242312
rect 405702 242256 408204 242312
rect 405641 242254 408204 242256
rect 434621 242312 436172 242314
rect 434621 242256 434626 242312
rect 434682 242256 436172 242312
rect 434621 242254 436172 242256
rect 462221 242312 464140 242314
rect 462221 242256 462226 242312
rect 462282 242256 464140 242312
rect 462221 242254 464140 242256
rect 489821 242312 492108 242314
rect 489821 242256 489826 242312
rect 489882 242256 492108 242312
rect 489821 242254 492108 242256
rect 518801 242312 520076 242314
rect 518801 242256 518806 242312
rect 518862 242256 520076 242312
rect 518801 242254 520076 242256
rect 545757 242312 548044 242314
rect 545757 242256 545762 242312
rect 545818 242256 548044 242312
rect 545757 242254 548044 242256
rect 13721 242251 13787 242254
rect 42701 242251 42767 242254
rect 70301 242251 70367 242254
rect 97901 242251 97967 242254
rect 126881 242251 126947 242254
rect 154481 242251 154547 242254
rect 182081 242251 182147 242254
rect 209681 242251 209747 242254
rect 238661 242251 238727 242254
rect 266261 242251 266327 242254
rect 293861 242251 293927 242254
rect 322841 242251 322907 242254
rect 350441 242251 350507 242254
rect 378041 242251 378107 242254
rect 405641 242251 405707 242254
rect 434621 242251 434687 242254
rect 462221 242251 462287 242254
rect 489821 242251 489887 242254
rect 518801 242251 518867 242254
rect 545757 242251 545823 242254
rect 37917 241634 37983 241637
rect 66253 241634 66319 241637
rect 93853 241634 93919 241637
rect 121453 241634 121519 241637
rect 149053 241634 149119 241637
rect 178033 241634 178099 241637
rect 205633 241634 205699 241637
rect 233233 241634 233299 241637
rect 262213 241634 262279 241637
rect 289813 241634 289879 241637
rect 317413 241634 317479 241637
rect 345013 241634 345079 241637
rect 373993 241634 374059 241637
rect 401593 241634 401659 241637
rect 429193 241634 429259 241637
rect 458173 241634 458239 241637
rect 485773 241634 485839 241637
rect 513373 241634 513439 241637
rect 542353 241634 542419 241637
rect 569953 241634 570019 241637
rect 35788 241632 37983 241634
rect 35788 241576 37922 241632
rect 37978 241576 37983 241632
rect 35788 241574 37983 241576
rect 63940 241632 66319 241634
rect 63940 241576 66258 241632
rect 66314 241576 66319 241632
rect 63940 241574 66319 241576
rect 91908 241632 93919 241634
rect 91908 241576 93858 241632
rect 93914 241576 93919 241632
rect 91908 241574 93919 241576
rect 119876 241632 121519 241634
rect 119876 241576 121458 241632
rect 121514 241576 121519 241632
rect 119876 241574 121519 241576
rect 147844 241632 149119 241634
rect 147844 241576 149058 241632
rect 149114 241576 149119 241632
rect 147844 241574 149119 241576
rect 175812 241632 178099 241634
rect 175812 241576 178038 241632
rect 178094 241576 178099 241632
rect 175812 241574 178099 241576
rect 203964 241632 205699 241634
rect 203964 241576 205638 241632
rect 205694 241576 205699 241632
rect 203964 241574 205699 241576
rect 231932 241632 233299 241634
rect 231932 241576 233238 241632
rect 233294 241576 233299 241632
rect 231932 241574 233299 241576
rect 259900 241632 262279 241634
rect 259900 241576 262218 241632
rect 262274 241576 262279 241632
rect 259900 241574 262279 241576
rect 287868 241632 289879 241634
rect 287868 241576 289818 241632
rect 289874 241576 289879 241632
rect 287868 241574 289879 241576
rect 315836 241632 317479 241634
rect 315836 241576 317418 241632
rect 317474 241576 317479 241632
rect 315836 241574 317479 241576
rect 343804 241632 345079 241634
rect 343804 241576 345018 241632
rect 345074 241576 345079 241632
rect 343804 241574 345079 241576
rect 371956 241632 374059 241634
rect 371956 241576 373998 241632
rect 374054 241576 374059 241632
rect 371956 241574 374059 241576
rect 399924 241632 401659 241634
rect 399924 241576 401598 241632
rect 401654 241576 401659 241632
rect 399924 241574 401659 241576
rect 427892 241632 429259 241634
rect 427892 241576 429198 241632
rect 429254 241576 429259 241632
rect 427892 241574 429259 241576
rect 455860 241632 458239 241634
rect 455860 241576 458178 241632
rect 458234 241576 458239 241632
rect 455860 241574 458239 241576
rect 483828 241632 485839 241634
rect 483828 241576 485778 241632
rect 485834 241576 485839 241632
rect 483828 241574 485839 241576
rect 511796 241632 513439 241634
rect 511796 241576 513378 241632
rect 513434 241576 513439 241632
rect 511796 241574 513439 241576
rect 539948 241632 542419 241634
rect 539948 241576 542358 241632
rect 542414 241576 542419 241632
rect 539948 241574 542419 241576
rect 567916 241632 570019 241634
rect 567916 241576 569958 241632
rect 570014 241576 570019 241632
rect 567916 241574 570019 241576
rect 37917 241571 37983 241574
rect 66253 241571 66319 241574
rect 93853 241571 93919 241574
rect 121453 241571 121519 241574
rect 149053 241571 149119 241574
rect 178033 241571 178099 241574
rect 205633 241571 205699 241574
rect 233233 241571 233299 241574
rect 262213 241571 262279 241574
rect 289813 241571 289879 241574
rect 317413 241571 317479 241574
rect 345013 241571 345079 241574
rect 373993 241571 374059 241574
rect 401593 241571 401659 241574
rect 429193 241571 429259 241574
rect 458173 241571 458239 241574
rect 485773 241571 485839 241574
rect 513373 241571 513439 241574
rect 542353 241571 542419 241574
rect 569953 241571 570019 241574
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect 13721 215250 13787 215253
rect 42701 215250 42767 215253
rect 97901 215250 97967 215253
rect 126881 215250 126947 215253
rect 154481 215250 154547 215253
rect 182081 215250 182147 215253
rect 209681 215250 209747 215253
rect 238661 215250 238727 215253
rect 266261 215250 266327 215253
rect 293861 215250 293927 215253
rect 322841 215250 322907 215253
rect 350441 215250 350507 215253
rect 378041 215250 378107 215253
rect 405641 215250 405707 215253
rect 434621 215250 434687 215253
rect 462221 215250 462287 215253
rect 489821 215250 489887 215253
rect 518801 215250 518867 215253
rect 545757 215250 545823 215253
rect 13721 215248 16100 215250
rect 13721 215192 13726 215248
rect 13782 215192 16100 215248
rect 13721 215190 16100 215192
rect 42701 215248 44068 215250
rect 42701 215192 42706 215248
rect 42762 215192 44068 215248
rect 97901 215248 100188 215250
rect 42701 215190 44068 215192
rect 13721 215187 13787 215190
rect 42701 215187 42767 215190
rect -960 214828 480 215068
rect 70301 214706 70367 214709
rect 72006 214706 72066 215220
rect 97901 215192 97906 215248
rect 97962 215192 100188 215248
rect 97901 215190 100188 215192
rect 126881 215248 128156 215250
rect 126881 215192 126886 215248
rect 126942 215192 128156 215248
rect 126881 215190 128156 215192
rect 154481 215248 156124 215250
rect 154481 215192 154486 215248
rect 154542 215192 156124 215248
rect 154481 215190 156124 215192
rect 182081 215248 184092 215250
rect 182081 215192 182086 215248
rect 182142 215192 184092 215248
rect 182081 215190 184092 215192
rect 209681 215248 212060 215250
rect 209681 215192 209686 215248
rect 209742 215192 212060 215248
rect 209681 215190 212060 215192
rect 238661 215248 240212 215250
rect 238661 215192 238666 215248
rect 238722 215192 240212 215248
rect 238661 215190 240212 215192
rect 266261 215248 268180 215250
rect 266261 215192 266266 215248
rect 266322 215192 268180 215248
rect 266261 215190 268180 215192
rect 293861 215248 296148 215250
rect 293861 215192 293866 215248
rect 293922 215192 296148 215248
rect 293861 215190 296148 215192
rect 322841 215248 324116 215250
rect 322841 215192 322846 215248
rect 322902 215192 324116 215248
rect 322841 215190 324116 215192
rect 350441 215248 352084 215250
rect 350441 215192 350446 215248
rect 350502 215192 352084 215248
rect 350441 215190 352084 215192
rect 378041 215248 380052 215250
rect 378041 215192 378046 215248
rect 378102 215192 380052 215248
rect 378041 215190 380052 215192
rect 405641 215248 408204 215250
rect 405641 215192 405646 215248
rect 405702 215192 408204 215248
rect 405641 215190 408204 215192
rect 434621 215248 436172 215250
rect 434621 215192 434626 215248
rect 434682 215192 436172 215248
rect 434621 215190 436172 215192
rect 462221 215248 464140 215250
rect 462221 215192 462226 215248
rect 462282 215192 464140 215248
rect 462221 215190 464140 215192
rect 489821 215248 492108 215250
rect 489821 215192 489826 215248
rect 489882 215192 492108 215248
rect 489821 215190 492108 215192
rect 518801 215248 520076 215250
rect 518801 215192 518806 215248
rect 518862 215192 520076 215248
rect 518801 215190 520076 215192
rect 545757 215248 548044 215250
rect 545757 215192 545762 215248
rect 545818 215192 548044 215248
rect 545757 215190 548044 215192
rect 97901 215187 97967 215190
rect 126881 215187 126947 215190
rect 154481 215187 154547 215190
rect 182081 215187 182147 215190
rect 209681 215187 209747 215190
rect 238661 215187 238727 215190
rect 266261 215187 266327 215190
rect 293861 215187 293927 215190
rect 322841 215187 322907 215190
rect 350441 215187 350507 215190
rect 378041 215187 378107 215190
rect 405641 215187 405707 215190
rect 434621 215187 434687 215190
rect 462221 215187 462287 215190
rect 489821 215187 489887 215190
rect 518801 215187 518867 215190
rect 545757 215187 545823 215190
rect 70301 214704 72066 214706
rect 70301 214648 70306 214704
rect 70362 214648 72066 214704
rect 70301 214646 72066 214648
rect 70301 214643 70367 214646
rect 37917 214570 37983 214573
rect 66253 214570 66319 214573
rect 93853 214570 93919 214573
rect 121453 214570 121519 214573
rect 149053 214570 149119 214573
rect 178033 214570 178099 214573
rect 233233 214570 233299 214573
rect 262213 214570 262279 214573
rect 289813 214570 289879 214573
rect 317413 214570 317479 214573
rect 345013 214570 345079 214573
rect 373993 214570 374059 214573
rect 401593 214570 401659 214573
rect 429193 214570 429259 214573
rect 458173 214570 458239 214573
rect 485773 214570 485839 214573
rect 513373 214570 513439 214573
rect 542353 214570 542419 214573
rect 569953 214570 570019 214573
rect 35788 214568 37983 214570
rect 35788 214512 37922 214568
rect 37978 214512 37983 214568
rect 35788 214510 37983 214512
rect 63940 214568 66319 214570
rect 63940 214512 66258 214568
rect 66314 214512 66319 214568
rect 63940 214510 66319 214512
rect 91908 214568 93919 214570
rect 91908 214512 93858 214568
rect 93914 214512 93919 214568
rect 91908 214510 93919 214512
rect 119876 214568 121519 214570
rect 119876 214512 121458 214568
rect 121514 214512 121519 214568
rect 119876 214510 121519 214512
rect 147844 214568 149119 214570
rect 147844 214512 149058 214568
rect 149114 214512 149119 214568
rect 147844 214510 149119 214512
rect 175812 214568 178099 214570
rect 175812 214512 178038 214568
rect 178094 214512 178099 214568
rect 231932 214568 233299 214570
rect 175812 214510 178099 214512
rect 37917 214507 37983 214510
rect 66253 214507 66319 214510
rect 93853 214507 93919 214510
rect 121453 214507 121519 214510
rect 149053 214507 149119 214510
rect 178033 214507 178099 214510
rect 203934 214026 203994 214540
rect 231932 214512 233238 214568
rect 233294 214512 233299 214568
rect 231932 214510 233299 214512
rect 259900 214568 262279 214570
rect 259900 214512 262218 214568
rect 262274 214512 262279 214568
rect 259900 214510 262279 214512
rect 287868 214568 289879 214570
rect 287868 214512 289818 214568
rect 289874 214512 289879 214568
rect 287868 214510 289879 214512
rect 315836 214568 317479 214570
rect 315836 214512 317418 214568
rect 317474 214512 317479 214568
rect 315836 214510 317479 214512
rect 343804 214568 345079 214570
rect 343804 214512 345018 214568
rect 345074 214512 345079 214568
rect 343804 214510 345079 214512
rect 371956 214568 374059 214570
rect 371956 214512 373998 214568
rect 374054 214512 374059 214568
rect 371956 214510 374059 214512
rect 399924 214568 401659 214570
rect 399924 214512 401598 214568
rect 401654 214512 401659 214568
rect 399924 214510 401659 214512
rect 427892 214568 429259 214570
rect 427892 214512 429198 214568
rect 429254 214512 429259 214568
rect 427892 214510 429259 214512
rect 455860 214568 458239 214570
rect 455860 214512 458178 214568
rect 458234 214512 458239 214568
rect 455860 214510 458239 214512
rect 483828 214568 485839 214570
rect 483828 214512 485778 214568
rect 485834 214512 485839 214568
rect 483828 214510 485839 214512
rect 511796 214568 513439 214570
rect 511796 214512 513378 214568
rect 513434 214512 513439 214568
rect 511796 214510 513439 214512
rect 539948 214568 542419 214570
rect 539948 214512 542358 214568
rect 542414 214512 542419 214568
rect 539948 214510 542419 214512
rect 567916 214568 570019 214570
rect 567916 214512 569958 214568
rect 570014 214512 570019 214568
rect 567916 214510 570019 214512
rect 233233 214507 233299 214510
rect 262213 214507 262279 214510
rect 289813 214507 289879 214510
rect 317413 214507 317479 214510
rect 345013 214507 345079 214510
rect 373993 214507 374059 214510
rect 401593 214507 401659 214510
rect 429193 214507 429259 214510
rect 458173 214507 458239 214510
rect 485773 214507 485839 214510
rect 513373 214507 513439 214510
rect 542353 214507 542419 214510
rect 569953 214507 570019 214510
rect 205633 214026 205699 214029
rect 203934 214024 205699 214026
rect 203934 213968 205638 214024
rect 205694 213968 205699 214024
rect 203934 213966 205699 213968
rect 205633 213963 205699 213966
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3785 201922 3851 201925
rect -960 201920 3851 201922
rect -960 201864 3790 201920
rect 3846 201864 3851 201920
rect -960 201862 3851 201864
rect -960 201772 480 201862
rect 3785 201859 3851 201862
rect 583520 192388 584960 192628
rect -960 188866 480 188956
rect 2957 188866 3023 188869
rect -960 188864 3023 188866
rect -960 188808 2962 188864
rect 3018 188808 3023 188864
rect -960 188806 3023 188808
rect -960 188716 480 188806
rect 2957 188803 3023 188806
rect 13721 188322 13787 188325
rect 42701 188322 42767 188325
rect 70301 188322 70367 188325
rect 97901 188322 97967 188325
rect 126881 188322 126947 188325
rect 154481 188322 154547 188325
rect 182081 188322 182147 188325
rect 209681 188322 209747 188325
rect 238661 188322 238727 188325
rect 266261 188322 266327 188325
rect 293861 188322 293927 188325
rect 322841 188322 322907 188325
rect 350441 188322 350507 188325
rect 378041 188322 378107 188325
rect 405641 188322 405707 188325
rect 434621 188322 434687 188325
rect 462221 188322 462287 188325
rect 489821 188322 489887 188325
rect 518801 188322 518867 188325
rect 545757 188322 545823 188325
rect 13721 188320 16100 188322
rect 13721 188264 13726 188320
rect 13782 188264 16100 188320
rect 13721 188262 16100 188264
rect 42701 188320 44068 188322
rect 42701 188264 42706 188320
rect 42762 188264 44068 188320
rect 42701 188262 44068 188264
rect 70301 188320 72036 188322
rect 70301 188264 70306 188320
rect 70362 188264 72036 188320
rect 70301 188262 72036 188264
rect 97901 188320 100188 188322
rect 97901 188264 97906 188320
rect 97962 188264 100188 188320
rect 97901 188262 100188 188264
rect 126881 188320 128156 188322
rect 126881 188264 126886 188320
rect 126942 188264 128156 188320
rect 126881 188262 128156 188264
rect 154481 188320 156124 188322
rect 154481 188264 154486 188320
rect 154542 188264 156124 188320
rect 154481 188262 156124 188264
rect 182081 188320 184092 188322
rect 182081 188264 182086 188320
rect 182142 188264 184092 188320
rect 182081 188262 184092 188264
rect 209681 188320 212060 188322
rect 209681 188264 209686 188320
rect 209742 188264 212060 188320
rect 209681 188262 212060 188264
rect 238661 188320 240212 188322
rect 238661 188264 238666 188320
rect 238722 188264 240212 188320
rect 238661 188262 240212 188264
rect 266261 188320 268180 188322
rect 266261 188264 266266 188320
rect 266322 188264 268180 188320
rect 266261 188262 268180 188264
rect 293861 188320 296148 188322
rect 293861 188264 293866 188320
rect 293922 188264 296148 188320
rect 293861 188262 296148 188264
rect 322841 188320 324116 188322
rect 322841 188264 322846 188320
rect 322902 188264 324116 188320
rect 322841 188262 324116 188264
rect 350441 188320 352084 188322
rect 350441 188264 350446 188320
rect 350502 188264 352084 188320
rect 350441 188262 352084 188264
rect 378041 188320 380052 188322
rect 378041 188264 378046 188320
rect 378102 188264 380052 188320
rect 378041 188262 380052 188264
rect 405641 188320 408204 188322
rect 405641 188264 405646 188320
rect 405702 188264 408204 188320
rect 405641 188262 408204 188264
rect 434621 188320 436172 188322
rect 434621 188264 434626 188320
rect 434682 188264 436172 188320
rect 434621 188262 436172 188264
rect 462221 188320 464140 188322
rect 462221 188264 462226 188320
rect 462282 188264 464140 188320
rect 462221 188262 464140 188264
rect 489821 188320 492108 188322
rect 489821 188264 489826 188320
rect 489882 188264 492108 188320
rect 489821 188262 492108 188264
rect 518801 188320 520076 188322
rect 518801 188264 518806 188320
rect 518862 188264 520076 188320
rect 518801 188262 520076 188264
rect 545757 188320 548044 188322
rect 545757 188264 545762 188320
rect 545818 188264 548044 188320
rect 545757 188262 548044 188264
rect 13721 188259 13787 188262
rect 42701 188259 42767 188262
rect 70301 188259 70367 188262
rect 97901 188259 97967 188262
rect 126881 188259 126947 188262
rect 154481 188259 154547 188262
rect 182081 188259 182147 188262
rect 209681 188259 209747 188262
rect 238661 188259 238727 188262
rect 266261 188259 266327 188262
rect 293861 188259 293927 188262
rect 322841 188259 322907 188262
rect 350441 188259 350507 188262
rect 378041 188259 378107 188262
rect 405641 188259 405707 188262
rect 434621 188259 434687 188262
rect 462221 188259 462287 188262
rect 489821 188259 489887 188262
rect 518801 188259 518867 188262
rect 545757 188259 545823 188262
rect 37917 187642 37983 187645
rect 66253 187642 66319 187645
rect 93853 187642 93919 187645
rect 121453 187642 121519 187645
rect 149053 187642 149119 187645
rect 178033 187642 178099 187645
rect 205633 187642 205699 187645
rect 233233 187642 233299 187645
rect 262213 187642 262279 187645
rect 289813 187642 289879 187645
rect 317413 187642 317479 187645
rect 345013 187642 345079 187645
rect 373993 187642 374059 187645
rect 401593 187642 401659 187645
rect 429193 187642 429259 187645
rect 458173 187642 458239 187645
rect 485773 187642 485839 187645
rect 513373 187642 513439 187645
rect 542353 187642 542419 187645
rect 569953 187642 570019 187645
rect 35788 187640 37983 187642
rect 35788 187584 37922 187640
rect 37978 187584 37983 187640
rect 35788 187582 37983 187584
rect 63940 187640 66319 187642
rect 63940 187584 66258 187640
rect 66314 187584 66319 187640
rect 63940 187582 66319 187584
rect 91908 187640 93919 187642
rect 91908 187584 93858 187640
rect 93914 187584 93919 187640
rect 91908 187582 93919 187584
rect 119876 187640 121519 187642
rect 119876 187584 121458 187640
rect 121514 187584 121519 187640
rect 119876 187582 121519 187584
rect 147844 187640 149119 187642
rect 147844 187584 149058 187640
rect 149114 187584 149119 187640
rect 147844 187582 149119 187584
rect 175812 187640 178099 187642
rect 175812 187584 178038 187640
rect 178094 187584 178099 187640
rect 175812 187582 178099 187584
rect 203964 187640 205699 187642
rect 203964 187584 205638 187640
rect 205694 187584 205699 187640
rect 203964 187582 205699 187584
rect 231932 187640 233299 187642
rect 231932 187584 233238 187640
rect 233294 187584 233299 187640
rect 231932 187582 233299 187584
rect 259900 187640 262279 187642
rect 259900 187584 262218 187640
rect 262274 187584 262279 187640
rect 259900 187582 262279 187584
rect 287868 187640 289879 187642
rect 287868 187584 289818 187640
rect 289874 187584 289879 187640
rect 287868 187582 289879 187584
rect 315836 187640 317479 187642
rect 315836 187584 317418 187640
rect 317474 187584 317479 187640
rect 315836 187582 317479 187584
rect 343804 187640 345079 187642
rect 343804 187584 345018 187640
rect 345074 187584 345079 187640
rect 343804 187582 345079 187584
rect 371956 187640 374059 187642
rect 371956 187584 373998 187640
rect 374054 187584 374059 187640
rect 371956 187582 374059 187584
rect 399924 187640 401659 187642
rect 399924 187584 401598 187640
rect 401654 187584 401659 187640
rect 399924 187582 401659 187584
rect 427892 187640 429259 187642
rect 427892 187584 429198 187640
rect 429254 187584 429259 187640
rect 427892 187582 429259 187584
rect 455860 187640 458239 187642
rect 455860 187584 458178 187640
rect 458234 187584 458239 187640
rect 455860 187582 458239 187584
rect 483828 187640 485839 187642
rect 483828 187584 485778 187640
rect 485834 187584 485839 187640
rect 483828 187582 485839 187584
rect 511796 187640 513439 187642
rect 511796 187584 513378 187640
rect 513434 187584 513439 187640
rect 511796 187582 513439 187584
rect 539948 187640 542419 187642
rect 539948 187584 542358 187640
rect 542414 187584 542419 187640
rect 539948 187582 542419 187584
rect 567916 187640 570019 187642
rect 567916 187584 569958 187640
rect 570014 187584 570019 187640
rect 567916 187582 570019 187584
rect 37917 187579 37983 187582
rect 66253 187579 66319 187582
rect 93853 187579 93919 187582
rect 121453 187579 121519 187582
rect 149053 187579 149119 187582
rect 178033 187579 178099 187582
rect 205633 187579 205699 187582
rect 233233 187579 233299 187582
rect 262213 187579 262279 187582
rect 289813 187579 289879 187582
rect 317413 187579 317479 187582
rect 345013 187579 345079 187582
rect 373993 187579 374059 187582
rect 401593 187579 401659 187582
rect 429193 187579 429259 187582
rect 458173 187579 458239 187582
rect 485773 187579 485839 187582
rect 513373 187579 513439 187582
rect 542353 187579 542419 187582
rect 569953 187579 570019 187582
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 13721 161258 13787 161261
rect 42701 161258 42767 161261
rect 70301 161258 70367 161261
rect 97901 161258 97967 161261
rect 126881 161258 126947 161261
rect 154481 161258 154547 161261
rect 182081 161258 182147 161261
rect 209681 161258 209747 161261
rect 238661 161258 238727 161261
rect 266261 161258 266327 161261
rect 293861 161258 293927 161261
rect 322841 161258 322907 161261
rect 350441 161258 350507 161261
rect 378041 161258 378107 161261
rect 405641 161258 405707 161261
rect 434621 161258 434687 161261
rect 462221 161258 462287 161261
rect 489821 161258 489887 161261
rect 518801 161258 518867 161261
rect 545757 161258 545823 161261
rect 13721 161256 16100 161258
rect 13721 161200 13726 161256
rect 13782 161200 16100 161256
rect 13721 161198 16100 161200
rect 42701 161256 44068 161258
rect 42701 161200 42706 161256
rect 42762 161200 44068 161256
rect 42701 161198 44068 161200
rect 70301 161256 72036 161258
rect 70301 161200 70306 161256
rect 70362 161200 72036 161256
rect 70301 161198 72036 161200
rect 97901 161256 100188 161258
rect 97901 161200 97906 161256
rect 97962 161200 100188 161256
rect 97901 161198 100188 161200
rect 126881 161256 128156 161258
rect 126881 161200 126886 161256
rect 126942 161200 128156 161256
rect 126881 161198 128156 161200
rect 154481 161256 156124 161258
rect 154481 161200 154486 161256
rect 154542 161200 156124 161256
rect 154481 161198 156124 161200
rect 182081 161256 184092 161258
rect 182081 161200 182086 161256
rect 182142 161200 184092 161256
rect 182081 161198 184092 161200
rect 209681 161256 212060 161258
rect 209681 161200 209686 161256
rect 209742 161200 212060 161256
rect 209681 161198 212060 161200
rect 238661 161256 240212 161258
rect 238661 161200 238666 161256
rect 238722 161200 240212 161256
rect 238661 161198 240212 161200
rect 266261 161256 268180 161258
rect 266261 161200 266266 161256
rect 266322 161200 268180 161256
rect 266261 161198 268180 161200
rect 293861 161256 296148 161258
rect 293861 161200 293866 161256
rect 293922 161200 296148 161256
rect 293861 161198 296148 161200
rect 322841 161256 324116 161258
rect 322841 161200 322846 161256
rect 322902 161200 324116 161256
rect 322841 161198 324116 161200
rect 350441 161256 352084 161258
rect 350441 161200 350446 161256
rect 350502 161200 352084 161256
rect 350441 161198 352084 161200
rect 378041 161256 380052 161258
rect 378041 161200 378046 161256
rect 378102 161200 380052 161256
rect 378041 161198 380052 161200
rect 405641 161256 408204 161258
rect 405641 161200 405646 161256
rect 405702 161200 408204 161256
rect 405641 161198 408204 161200
rect 434621 161256 436172 161258
rect 434621 161200 434626 161256
rect 434682 161200 436172 161256
rect 434621 161198 436172 161200
rect 462221 161256 464140 161258
rect 462221 161200 462226 161256
rect 462282 161200 464140 161256
rect 462221 161198 464140 161200
rect 489821 161256 492108 161258
rect 489821 161200 489826 161256
rect 489882 161200 492108 161256
rect 489821 161198 492108 161200
rect 518801 161256 520076 161258
rect 518801 161200 518806 161256
rect 518862 161200 520076 161256
rect 518801 161198 520076 161200
rect 545757 161256 548044 161258
rect 545757 161200 545762 161256
rect 545818 161200 548044 161256
rect 545757 161198 548044 161200
rect 13721 161195 13787 161198
rect 42701 161195 42767 161198
rect 70301 161195 70367 161198
rect 97901 161195 97967 161198
rect 126881 161195 126947 161198
rect 154481 161195 154547 161198
rect 182081 161195 182147 161198
rect 209681 161195 209747 161198
rect 238661 161195 238727 161198
rect 266261 161195 266327 161198
rect 293861 161195 293927 161198
rect 322841 161195 322907 161198
rect 350441 161195 350507 161198
rect 378041 161195 378107 161198
rect 405641 161195 405707 161198
rect 434621 161195 434687 161198
rect 462221 161195 462287 161198
rect 489821 161195 489887 161198
rect 518801 161195 518867 161198
rect 545757 161195 545823 161198
rect 37917 160578 37983 160581
rect 66253 160578 66319 160581
rect 93853 160578 93919 160581
rect 121453 160578 121519 160581
rect 149053 160578 149119 160581
rect 178033 160578 178099 160581
rect 205633 160578 205699 160581
rect 233233 160578 233299 160581
rect 262213 160578 262279 160581
rect 289813 160578 289879 160581
rect 317413 160578 317479 160581
rect 345013 160578 345079 160581
rect 373993 160578 374059 160581
rect 401593 160578 401659 160581
rect 429193 160578 429259 160581
rect 458173 160578 458239 160581
rect 485773 160578 485839 160581
rect 513373 160578 513439 160581
rect 542353 160578 542419 160581
rect 569953 160578 570019 160581
rect 35788 160576 37983 160578
rect 35788 160520 37922 160576
rect 37978 160520 37983 160576
rect 35788 160518 37983 160520
rect 63940 160576 66319 160578
rect 63940 160520 66258 160576
rect 66314 160520 66319 160576
rect 63940 160518 66319 160520
rect 91908 160576 93919 160578
rect 91908 160520 93858 160576
rect 93914 160520 93919 160576
rect 91908 160518 93919 160520
rect 119876 160576 121519 160578
rect 119876 160520 121458 160576
rect 121514 160520 121519 160576
rect 119876 160518 121519 160520
rect 147844 160576 149119 160578
rect 147844 160520 149058 160576
rect 149114 160520 149119 160576
rect 147844 160518 149119 160520
rect 175812 160576 178099 160578
rect 175812 160520 178038 160576
rect 178094 160520 178099 160576
rect 175812 160518 178099 160520
rect 203964 160576 205699 160578
rect 203964 160520 205638 160576
rect 205694 160520 205699 160576
rect 203964 160518 205699 160520
rect 231932 160576 233299 160578
rect 231932 160520 233238 160576
rect 233294 160520 233299 160576
rect 231932 160518 233299 160520
rect 259900 160576 262279 160578
rect 259900 160520 262218 160576
rect 262274 160520 262279 160576
rect 259900 160518 262279 160520
rect 287868 160576 289879 160578
rect 287868 160520 289818 160576
rect 289874 160520 289879 160576
rect 287868 160518 289879 160520
rect 315836 160576 317479 160578
rect 315836 160520 317418 160576
rect 317474 160520 317479 160576
rect 315836 160518 317479 160520
rect 343804 160576 345079 160578
rect 343804 160520 345018 160576
rect 345074 160520 345079 160576
rect 343804 160518 345079 160520
rect 371956 160576 374059 160578
rect 371956 160520 373998 160576
rect 374054 160520 374059 160576
rect 371956 160518 374059 160520
rect 399924 160576 401659 160578
rect 399924 160520 401598 160576
rect 401654 160520 401659 160576
rect 399924 160518 401659 160520
rect 427892 160576 429259 160578
rect 427892 160520 429198 160576
rect 429254 160520 429259 160576
rect 427892 160518 429259 160520
rect 455860 160576 458239 160578
rect 455860 160520 458178 160576
rect 458234 160520 458239 160576
rect 455860 160518 458239 160520
rect 483828 160576 485839 160578
rect 483828 160520 485778 160576
rect 485834 160520 485839 160576
rect 483828 160518 485839 160520
rect 511796 160576 513439 160578
rect 511796 160520 513378 160576
rect 513434 160520 513439 160576
rect 511796 160518 513439 160520
rect 539948 160576 542419 160578
rect 539948 160520 542358 160576
rect 542414 160520 542419 160576
rect 539948 160518 542419 160520
rect 567916 160576 570019 160578
rect 567916 160520 569958 160576
rect 570014 160520 570019 160576
rect 567916 160518 570019 160520
rect 37917 160515 37983 160518
rect 66253 160515 66319 160518
rect 93853 160515 93919 160518
rect 121453 160515 121519 160518
rect 149053 160515 149119 160518
rect 178033 160515 178099 160518
rect 205633 160515 205699 160518
rect 233233 160515 233299 160518
rect 262213 160515 262279 160518
rect 289813 160515 289879 160518
rect 317413 160515 317479 160518
rect 345013 160515 345079 160518
rect 373993 160515 374059 160518
rect 401593 160515 401659 160518
rect 429193 160515 429259 160518
rect 458173 160515 458239 160518
rect 485773 160515 485839 160518
rect 513373 160515 513439 160518
rect 542353 160515 542419 160518
rect 569953 160515 570019 160518
rect 583520 152540 584960 152780
rect -960 149834 480 149924
rect 3877 149834 3943 149837
rect -960 149832 3943 149834
rect -960 149776 3882 149832
rect 3938 149776 3943 149832
rect -960 149774 3943 149776
rect -960 149684 480 149774
rect 3877 149771 3943 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3969 136778 4035 136781
rect -960 136776 4035 136778
rect -960 136720 3974 136776
rect 4030 136720 4035 136776
rect -960 136718 4035 136720
rect -960 136628 480 136718
rect 3969 136715 4035 136718
rect 13721 134330 13787 134333
rect 42701 134330 42767 134333
rect 70301 134330 70367 134333
rect 97901 134330 97967 134333
rect 126881 134330 126947 134333
rect 154481 134330 154547 134333
rect 182081 134330 182147 134333
rect 209681 134330 209747 134333
rect 238661 134330 238727 134333
rect 266261 134330 266327 134333
rect 293861 134330 293927 134333
rect 322841 134330 322907 134333
rect 350441 134330 350507 134333
rect 378041 134330 378107 134333
rect 405641 134330 405707 134333
rect 434621 134330 434687 134333
rect 462221 134330 462287 134333
rect 489821 134330 489887 134333
rect 518801 134330 518867 134333
rect 545757 134330 545823 134333
rect 13721 134328 16100 134330
rect 13721 134272 13726 134328
rect 13782 134272 16100 134328
rect 13721 134270 16100 134272
rect 42701 134328 44068 134330
rect 42701 134272 42706 134328
rect 42762 134272 44068 134328
rect 42701 134270 44068 134272
rect 70301 134328 72036 134330
rect 70301 134272 70306 134328
rect 70362 134272 72036 134328
rect 70301 134270 72036 134272
rect 97901 134328 100188 134330
rect 97901 134272 97906 134328
rect 97962 134272 100188 134328
rect 97901 134270 100188 134272
rect 126881 134328 128156 134330
rect 126881 134272 126886 134328
rect 126942 134272 128156 134328
rect 126881 134270 128156 134272
rect 154481 134328 156124 134330
rect 154481 134272 154486 134328
rect 154542 134272 156124 134328
rect 154481 134270 156124 134272
rect 182081 134328 184092 134330
rect 182081 134272 182086 134328
rect 182142 134272 184092 134328
rect 182081 134270 184092 134272
rect 209681 134328 212060 134330
rect 209681 134272 209686 134328
rect 209742 134272 212060 134328
rect 209681 134270 212060 134272
rect 238661 134328 240212 134330
rect 238661 134272 238666 134328
rect 238722 134272 240212 134328
rect 238661 134270 240212 134272
rect 266261 134328 268180 134330
rect 266261 134272 266266 134328
rect 266322 134272 268180 134328
rect 266261 134270 268180 134272
rect 293861 134328 296148 134330
rect 293861 134272 293866 134328
rect 293922 134272 296148 134328
rect 293861 134270 296148 134272
rect 322841 134328 324116 134330
rect 322841 134272 322846 134328
rect 322902 134272 324116 134328
rect 322841 134270 324116 134272
rect 350441 134328 352084 134330
rect 350441 134272 350446 134328
rect 350502 134272 352084 134328
rect 350441 134270 352084 134272
rect 378041 134328 380052 134330
rect 378041 134272 378046 134328
rect 378102 134272 380052 134328
rect 378041 134270 380052 134272
rect 405641 134328 408204 134330
rect 405641 134272 405646 134328
rect 405702 134272 408204 134328
rect 405641 134270 408204 134272
rect 434621 134328 436172 134330
rect 434621 134272 434626 134328
rect 434682 134272 436172 134328
rect 434621 134270 436172 134272
rect 462221 134328 464140 134330
rect 462221 134272 462226 134328
rect 462282 134272 464140 134328
rect 462221 134270 464140 134272
rect 489821 134328 492108 134330
rect 489821 134272 489826 134328
rect 489882 134272 492108 134328
rect 489821 134270 492108 134272
rect 518801 134328 520076 134330
rect 518801 134272 518806 134328
rect 518862 134272 520076 134328
rect 518801 134270 520076 134272
rect 545757 134328 548044 134330
rect 545757 134272 545762 134328
rect 545818 134272 548044 134328
rect 545757 134270 548044 134272
rect 13721 134267 13787 134270
rect 42701 134267 42767 134270
rect 70301 134267 70367 134270
rect 97901 134267 97967 134270
rect 126881 134267 126947 134270
rect 154481 134267 154547 134270
rect 182081 134267 182147 134270
rect 209681 134267 209747 134270
rect 238661 134267 238727 134270
rect 266261 134267 266327 134270
rect 293861 134267 293927 134270
rect 322841 134267 322907 134270
rect 350441 134267 350507 134270
rect 378041 134267 378107 134270
rect 405641 134267 405707 134270
rect 434621 134267 434687 134270
rect 462221 134267 462287 134270
rect 489821 134267 489887 134270
rect 518801 134267 518867 134270
rect 545757 134267 545823 134270
rect 37917 133650 37983 133653
rect 66253 133650 66319 133653
rect 93853 133650 93919 133653
rect 121453 133650 121519 133653
rect 149053 133650 149119 133653
rect 178033 133650 178099 133653
rect 205633 133650 205699 133653
rect 233233 133650 233299 133653
rect 262213 133650 262279 133653
rect 289813 133650 289879 133653
rect 317413 133650 317479 133653
rect 345013 133650 345079 133653
rect 373993 133650 374059 133653
rect 401593 133650 401659 133653
rect 429193 133650 429259 133653
rect 458173 133650 458239 133653
rect 485773 133650 485839 133653
rect 513373 133650 513439 133653
rect 542353 133650 542419 133653
rect 569953 133650 570019 133653
rect 35788 133648 37983 133650
rect 35788 133592 37922 133648
rect 37978 133592 37983 133648
rect 35788 133590 37983 133592
rect 63940 133648 66319 133650
rect 63940 133592 66258 133648
rect 66314 133592 66319 133648
rect 63940 133590 66319 133592
rect 91908 133648 93919 133650
rect 91908 133592 93858 133648
rect 93914 133592 93919 133648
rect 91908 133590 93919 133592
rect 119876 133648 121519 133650
rect 119876 133592 121458 133648
rect 121514 133592 121519 133648
rect 119876 133590 121519 133592
rect 147844 133648 149119 133650
rect 147844 133592 149058 133648
rect 149114 133592 149119 133648
rect 147844 133590 149119 133592
rect 175812 133648 178099 133650
rect 175812 133592 178038 133648
rect 178094 133592 178099 133648
rect 175812 133590 178099 133592
rect 203964 133648 205699 133650
rect 203964 133592 205638 133648
rect 205694 133592 205699 133648
rect 203964 133590 205699 133592
rect 231932 133648 233299 133650
rect 231932 133592 233238 133648
rect 233294 133592 233299 133648
rect 231932 133590 233299 133592
rect 259900 133648 262279 133650
rect 259900 133592 262218 133648
rect 262274 133592 262279 133648
rect 259900 133590 262279 133592
rect 287868 133648 289879 133650
rect 287868 133592 289818 133648
rect 289874 133592 289879 133648
rect 287868 133590 289879 133592
rect 315836 133648 317479 133650
rect 315836 133592 317418 133648
rect 317474 133592 317479 133648
rect 315836 133590 317479 133592
rect 343804 133648 345079 133650
rect 343804 133592 345018 133648
rect 345074 133592 345079 133648
rect 343804 133590 345079 133592
rect 371956 133648 374059 133650
rect 371956 133592 373998 133648
rect 374054 133592 374059 133648
rect 371956 133590 374059 133592
rect 399924 133648 401659 133650
rect 399924 133592 401598 133648
rect 401654 133592 401659 133648
rect 399924 133590 401659 133592
rect 427892 133648 429259 133650
rect 427892 133592 429198 133648
rect 429254 133592 429259 133648
rect 427892 133590 429259 133592
rect 455860 133648 458239 133650
rect 455860 133592 458178 133648
rect 458234 133592 458239 133648
rect 455860 133590 458239 133592
rect 483828 133648 485839 133650
rect 483828 133592 485778 133648
rect 485834 133592 485839 133648
rect 483828 133590 485839 133592
rect 511796 133648 513439 133650
rect 511796 133592 513378 133648
rect 513434 133592 513439 133648
rect 511796 133590 513439 133592
rect 539948 133648 542419 133650
rect 539948 133592 542358 133648
rect 542414 133592 542419 133648
rect 539948 133590 542419 133592
rect 567916 133648 570019 133650
rect 567916 133592 569958 133648
rect 570014 133592 570019 133648
rect 567916 133590 570019 133592
rect 37917 133587 37983 133590
rect 66253 133587 66319 133590
rect 93853 133587 93919 133590
rect 121453 133587 121519 133590
rect 149053 133587 149119 133590
rect 178033 133587 178099 133590
rect 205633 133587 205699 133590
rect 233233 133587 233299 133590
rect 262213 133587 262279 133590
rect 289813 133587 289879 133590
rect 317413 133587 317479 133590
rect 345013 133587 345079 133590
rect 373993 133587 374059 133590
rect 401593 133587 401659 133590
rect 429193 133587 429259 133590
rect 458173 133587 458239 133590
rect 485773 133587 485839 133590
rect 513373 133587 513439 133590
rect 542353 133587 542419 133590
rect 569953 133587 570019 133590
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 13721 107266 13787 107269
rect 42701 107266 42767 107269
rect 70301 107266 70367 107269
rect 97901 107266 97967 107269
rect 126881 107266 126947 107269
rect 154481 107266 154547 107269
rect 182081 107266 182147 107269
rect 209681 107266 209747 107269
rect 238661 107266 238727 107269
rect 266261 107266 266327 107269
rect 293861 107266 293927 107269
rect 322841 107266 322907 107269
rect 350441 107266 350507 107269
rect 378041 107266 378107 107269
rect 405641 107266 405707 107269
rect 434621 107266 434687 107269
rect 462221 107266 462287 107269
rect 489821 107266 489887 107269
rect 518801 107266 518867 107269
rect 545757 107266 545823 107269
rect 13721 107264 16100 107266
rect 13721 107208 13726 107264
rect 13782 107208 16100 107264
rect 13721 107206 16100 107208
rect 42701 107264 44068 107266
rect 42701 107208 42706 107264
rect 42762 107208 44068 107264
rect 42701 107206 44068 107208
rect 70301 107264 72036 107266
rect 70301 107208 70306 107264
rect 70362 107208 72036 107264
rect 70301 107206 72036 107208
rect 97901 107264 100188 107266
rect 97901 107208 97906 107264
rect 97962 107208 100188 107264
rect 97901 107206 100188 107208
rect 126881 107264 128156 107266
rect 126881 107208 126886 107264
rect 126942 107208 128156 107264
rect 126881 107206 128156 107208
rect 154481 107264 156124 107266
rect 154481 107208 154486 107264
rect 154542 107208 156124 107264
rect 154481 107206 156124 107208
rect 182081 107264 184092 107266
rect 182081 107208 182086 107264
rect 182142 107208 184092 107264
rect 182081 107206 184092 107208
rect 209681 107264 212060 107266
rect 209681 107208 209686 107264
rect 209742 107208 212060 107264
rect 209681 107206 212060 107208
rect 238661 107264 240212 107266
rect 238661 107208 238666 107264
rect 238722 107208 240212 107264
rect 238661 107206 240212 107208
rect 266261 107264 268180 107266
rect 266261 107208 266266 107264
rect 266322 107208 268180 107264
rect 266261 107206 268180 107208
rect 293861 107264 296148 107266
rect 293861 107208 293866 107264
rect 293922 107208 296148 107264
rect 293861 107206 296148 107208
rect 322841 107264 324116 107266
rect 322841 107208 322846 107264
rect 322902 107208 324116 107264
rect 322841 107206 324116 107208
rect 350441 107264 352084 107266
rect 350441 107208 350446 107264
rect 350502 107208 352084 107264
rect 350441 107206 352084 107208
rect 378041 107264 380052 107266
rect 378041 107208 378046 107264
rect 378102 107208 380052 107264
rect 378041 107206 380052 107208
rect 405641 107264 408204 107266
rect 405641 107208 405646 107264
rect 405702 107208 408204 107264
rect 405641 107206 408204 107208
rect 434621 107264 436172 107266
rect 434621 107208 434626 107264
rect 434682 107208 436172 107264
rect 434621 107206 436172 107208
rect 462221 107264 464140 107266
rect 462221 107208 462226 107264
rect 462282 107208 464140 107264
rect 462221 107206 464140 107208
rect 489821 107264 492108 107266
rect 489821 107208 489826 107264
rect 489882 107208 492108 107264
rect 489821 107206 492108 107208
rect 518801 107264 520076 107266
rect 518801 107208 518806 107264
rect 518862 107208 520076 107264
rect 518801 107206 520076 107208
rect 545757 107264 548044 107266
rect 545757 107208 545762 107264
rect 545818 107208 548044 107264
rect 545757 107206 548044 107208
rect 13721 107203 13787 107206
rect 42701 107203 42767 107206
rect 70301 107203 70367 107206
rect 97901 107203 97967 107206
rect 126881 107203 126947 107206
rect 154481 107203 154547 107206
rect 182081 107203 182147 107206
rect 209681 107203 209747 107206
rect 238661 107203 238727 107206
rect 266261 107203 266327 107206
rect 293861 107203 293927 107206
rect 322841 107203 322907 107206
rect 350441 107203 350507 107206
rect 378041 107203 378107 107206
rect 405641 107203 405707 107206
rect 434621 107203 434687 107206
rect 462221 107203 462287 107206
rect 489821 107203 489887 107206
rect 518801 107203 518867 107206
rect 545757 107203 545823 107206
rect 37917 106586 37983 106589
rect 66253 106586 66319 106589
rect 93853 106586 93919 106589
rect 121453 106586 121519 106589
rect 149053 106586 149119 106589
rect 178033 106586 178099 106589
rect 205633 106586 205699 106589
rect 233233 106586 233299 106589
rect 262213 106586 262279 106589
rect 289813 106586 289879 106589
rect 317413 106586 317479 106589
rect 345013 106586 345079 106589
rect 373993 106586 374059 106589
rect 401593 106586 401659 106589
rect 429193 106586 429259 106589
rect 458173 106586 458239 106589
rect 485773 106586 485839 106589
rect 513373 106586 513439 106589
rect 542353 106586 542419 106589
rect 569953 106586 570019 106589
rect 35788 106584 37983 106586
rect 35788 106528 37922 106584
rect 37978 106528 37983 106584
rect 35788 106526 37983 106528
rect 63940 106584 66319 106586
rect 63940 106528 66258 106584
rect 66314 106528 66319 106584
rect 63940 106526 66319 106528
rect 91908 106584 93919 106586
rect 91908 106528 93858 106584
rect 93914 106528 93919 106584
rect 91908 106526 93919 106528
rect 119876 106584 121519 106586
rect 119876 106528 121458 106584
rect 121514 106528 121519 106584
rect 119876 106526 121519 106528
rect 147844 106584 149119 106586
rect 147844 106528 149058 106584
rect 149114 106528 149119 106584
rect 147844 106526 149119 106528
rect 175812 106584 178099 106586
rect 175812 106528 178038 106584
rect 178094 106528 178099 106584
rect 175812 106526 178099 106528
rect 203964 106584 205699 106586
rect 203964 106528 205638 106584
rect 205694 106528 205699 106584
rect 203964 106526 205699 106528
rect 231932 106584 233299 106586
rect 231932 106528 233238 106584
rect 233294 106528 233299 106584
rect 231932 106526 233299 106528
rect 259900 106584 262279 106586
rect 259900 106528 262218 106584
rect 262274 106528 262279 106584
rect 259900 106526 262279 106528
rect 287868 106584 289879 106586
rect 287868 106528 289818 106584
rect 289874 106528 289879 106584
rect 287868 106526 289879 106528
rect 315836 106584 317479 106586
rect 315836 106528 317418 106584
rect 317474 106528 317479 106584
rect 315836 106526 317479 106528
rect 343804 106584 345079 106586
rect 343804 106528 345018 106584
rect 345074 106528 345079 106584
rect 343804 106526 345079 106528
rect 371956 106584 374059 106586
rect 371956 106528 373998 106584
rect 374054 106528 374059 106584
rect 371956 106526 374059 106528
rect 399924 106584 401659 106586
rect 399924 106528 401598 106584
rect 401654 106528 401659 106584
rect 399924 106526 401659 106528
rect 427892 106584 429259 106586
rect 427892 106528 429198 106584
rect 429254 106528 429259 106584
rect 427892 106526 429259 106528
rect 455860 106584 458239 106586
rect 455860 106528 458178 106584
rect 458234 106528 458239 106584
rect 455860 106526 458239 106528
rect 483828 106584 485839 106586
rect 483828 106528 485778 106584
rect 485834 106528 485839 106584
rect 483828 106526 485839 106528
rect 511796 106584 513439 106586
rect 511796 106528 513378 106584
rect 513434 106528 513439 106584
rect 511796 106526 513439 106528
rect 539948 106584 542419 106586
rect 539948 106528 542358 106584
rect 542414 106528 542419 106584
rect 539948 106526 542419 106528
rect 567916 106584 570019 106586
rect 567916 106528 569958 106584
rect 570014 106528 570019 106584
rect 567916 106526 570019 106528
rect 37917 106523 37983 106526
rect 66253 106523 66319 106526
rect 93853 106523 93919 106526
rect 121453 106523 121519 106526
rect 149053 106523 149119 106526
rect 178033 106523 178099 106526
rect 205633 106523 205699 106526
rect 233233 106523 233299 106526
rect 262213 106523 262279 106526
rect 289813 106523 289879 106526
rect 317413 106523 317479 106526
rect 345013 106523 345079 106526
rect 373993 106523 374059 106526
rect 401593 106523 401659 106526
rect 429193 106523 429259 106526
rect 458173 106523 458239 106526
rect 485773 106523 485839 106526
rect 513373 106523 513439 106526
rect 542353 106523 542419 106526
rect 569953 106523 570019 106526
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 4061 97610 4127 97613
rect -960 97608 4127 97610
rect -960 97552 4066 97608
rect 4122 97552 4127 97608
rect -960 97550 4127 97552
rect -960 97460 480 97550
rect 4061 97547 4127 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 13721 80338 13787 80341
rect 42701 80338 42767 80341
rect 70301 80338 70367 80341
rect 97901 80338 97967 80341
rect 126881 80338 126947 80341
rect 154481 80338 154547 80341
rect 182081 80338 182147 80341
rect 209681 80338 209747 80341
rect 238661 80338 238727 80341
rect 266261 80338 266327 80341
rect 293861 80338 293927 80341
rect 322841 80338 322907 80341
rect 350441 80338 350507 80341
rect 378041 80338 378107 80341
rect 405641 80338 405707 80341
rect 434621 80338 434687 80341
rect 462221 80338 462287 80341
rect 489821 80338 489887 80341
rect 518801 80338 518867 80341
rect 545757 80338 545823 80341
rect 13721 80336 16100 80338
rect 13721 80280 13726 80336
rect 13782 80280 16100 80336
rect 13721 80278 16100 80280
rect 42701 80336 44068 80338
rect 42701 80280 42706 80336
rect 42762 80280 44068 80336
rect 42701 80278 44068 80280
rect 70301 80336 72036 80338
rect 70301 80280 70306 80336
rect 70362 80280 72036 80336
rect 70301 80278 72036 80280
rect 97901 80336 100188 80338
rect 97901 80280 97906 80336
rect 97962 80280 100188 80336
rect 97901 80278 100188 80280
rect 126881 80336 128156 80338
rect 126881 80280 126886 80336
rect 126942 80280 128156 80336
rect 126881 80278 128156 80280
rect 154481 80336 156124 80338
rect 154481 80280 154486 80336
rect 154542 80280 156124 80336
rect 154481 80278 156124 80280
rect 182081 80336 184092 80338
rect 182081 80280 182086 80336
rect 182142 80280 184092 80336
rect 182081 80278 184092 80280
rect 209681 80336 212060 80338
rect 209681 80280 209686 80336
rect 209742 80280 212060 80336
rect 209681 80278 212060 80280
rect 238661 80336 240212 80338
rect 238661 80280 238666 80336
rect 238722 80280 240212 80336
rect 238661 80278 240212 80280
rect 266261 80336 268180 80338
rect 266261 80280 266266 80336
rect 266322 80280 268180 80336
rect 266261 80278 268180 80280
rect 293861 80336 296148 80338
rect 293861 80280 293866 80336
rect 293922 80280 296148 80336
rect 293861 80278 296148 80280
rect 322841 80336 324116 80338
rect 322841 80280 322846 80336
rect 322902 80280 324116 80336
rect 322841 80278 324116 80280
rect 350441 80336 352084 80338
rect 350441 80280 350446 80336
rect 350502 80280 352084 80336
rect 350441 80278 352084 80280
rect 378041 80336 380052 80338
rect 378041 80280 378046 80336
rect 378102 80280 380052 80336
rect 378041 80278 380052 80280
rect 405641 80336 408204 80338
rect 405641 80280 405646 80336
rect 405702 80280 408204 80336
rect 405641 80278 408204 80280
rect 434621 80336 436172 80338
rect 434621 80280 434626 80336
rect 434682 80280 436172 80336
rect 434621 80278 436172 80280
rect 462221 80336 464140 80338
rect 462221 80280 462226 80336
rect 462282 80280 464140 80336
rect 462221 80278 464140 80280
rect 489821 80336 492108 80338
rect 489821 80280 489826 80336
rect 489882 80280 492108 80336
rect 489821 80278 492108 80280
rect 518801 80336 520076 80338
rect 518801 80280 518806 80336
rect 518862 80280 520076 80336
rect 518801 80278 520076 80280
rect 545757 80336 548044 80338
rect 545757 80280 545762 80336
rect 545818 80280 548044 80336
rect 545757 80278 548044 80280
rect 13721 80275 13787 80278
rect 42701 80275 42767 80278
rect 70301 80275 70367 80278
rect 97901 80275 97967 80278
rect 126881 80275 126947 80278
rect 154481 80275 154547 80278
rect 182081 80275 182147 80278
rect 209681 80275 209747 80278
rect 238661 80275 238727 80278
rect 266261 80275 266327 80278
rect 293861 80275 293927 80278
rect 322841 80275 322907 80278
rect 350441 80275 350507 80278
rect 378041 80275 378107 80278
rect 405641 80275 405707 80278
rect 434621 80275 434687 80278
rect 462221 80275 462287 80278
rect 489821 80275 489887 80278
rect 518801 80275 518867 80278
rect 545757 80275 545823 80278
rect 37917 79658 37983 79661
rect 66253 79658 66319 79661
rect 93853 79658 93919 79661
rect 121453 79658 121519 79661
rect 149053 79658 149119 79661
rect 178033 79658 178099 79661
rect 205633 79658 205699 79661
rect 233233 79658 233299 79661
rect 262213 79658 262279 79661
rect 289813 79658 289879 79661
rect 317413 79658 317479 79661
rect 345013 79658 345079 79661
rect 373993 79658 374059 79661
rect 401593 79658 401659 79661
rect 429193 79658 429259 79661
rect 458173 79658 458239 79661
rect 485773 79658 485839 79661
rect 513373 79658 513439 79661
rect 542353 79658 542419 79661
rect 569953 79658 570019 79661
rect 35788 79656 37983 79658
rect 35788 79600 37922 79656
rect 37978 79600 37983 79656
rect 35788 79598 37983 79600
rect 63940 79656 66319 79658
rect 63940 79600 66258 79656
rect 66314 79600 66319 79656
rect 63940 79598 66319 79600
rect 91908 79656 93919 79658
rect 91908 79600 93858 79656
rect 93914 79600 93919 79656
rect 91908 79598 93919 79600
rect 119876 79656 121519 79658
rect 119876 79600 121458 79656
rect 121514 79600 121519 79656
rect 119876 79598 121519 79600
rect 147844 79656 149119 79658
rect 147844 79600 149058 79656
rect 149114 79600 149119 79656
rect 147844 79598 149119 79600
rect 175812 79656 178099 79658
rect 175812 79600 178038 79656
rect 178094 79600 178099 79656
rect 175812 79598 178099 79600
rect 203964 79656 205699 79658
rect 203964 79600 205638 79656
rect 205694 79600 205699 79656
rect 203964 79598 205699 79600
rect 231932 79656 233299 79658
rect 231932 79600 233238 79656
rect 233294 79600 233299 79656
rect 231932 79598 233299 79600
rect 259900 79656 262279 79658
rect 259900 79600 262218 79656
rect 262274 79600 262279 79656
rect 259900 79598 262279 79600
rect 287868 79656 289879 79658
rect 287868 79600 289818 79656
rect 289874 79600 289879 79656
rect 287868 79598 289879 79600
rect 315836 79656 317479 79658
rect 315836 79600 317418 79656
rect 317474 79600 317479 79656
rect 315836 79598 317479 79600
rect 343804 79656 345079 79658
rect 343804 79600 345018 79656
rect 345074 79600 345079 79656
rect 343804 79598 345079 79600
rect 371956 79656 374059 79658
rect 371956 79600 373998 79656
rect 374054 79600 374059 79656
rect 371956 79598 374059 79600
rect 399924 79656 401659 79658
rect 399924 79600 401598 79656
rect 401654 79600 401659 79656
rect 399924 79598 401659 79600
rect 427892 79656 429259 79658
rect 427892 79600 429198 79656
rect 429254 79600 429259 79656
rect 427892 79598 429259 79600
rect 455860 79656 458239 79658
rect 455860 79600 458178 79656
rect 458234 79600 458239 79656
rect 455860 79598 458239 79600
rect 483828 79656 485839 79658
rect 483828 79600 485778 79656
rect 485834 79600 485839 79656
rect 483828 79598 485839 79600
rect 511796 79656 513439 79658
rect 511796 79600 513378 79656
rect 513434 79600 513439 79656
rect 511796 79598 513439 79600
rect 539948 79656 542419 79658
rect 539948 79600 542358 79656
rect 542414 79600 542419 79656
rect 539948 79598 542419 79600
rect 567916 79656 570019 79658
rect 567916 79600 569958 79656
rect 570014 79600 570019 79656
rect 567916 79598 570019 79600
rect 37917 79595 37983 79598
rect 66253 79595 66319 79598
rect 93853 79595 93919 79598
rect 121453 79595 121519 79598
rect 149053 79595 149119 79598
rect 178033 79595 178099 79598
rect 205633 79595 205699 79598
rect 233233 79595 233299 79598
rect 262213 79595 262279 79598
rect 289813 79595 289879 79598
rect 317413 79595 317479 79598
rect 345013 79595 345079 79598
rect 373993 79595 374059 79598
rect 401593 79595 401659 79598
rect 429193 79595 429259 79598
rect 458173 79595 458239 79598
rect 485773 79595 485839 79598
rect 513373 79595 513439 79598
rect 542353 79595 542419 79598
rect 569953 79595 570019 79598
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 13721 53274 13787 53277
rect 42701 53274 42767 53277
rect 70301 53274 70367 53277
rect 97901 53274 97967 53277
rect 126881 53274 126947 53277
rect 154481 53274 154547 53277
rect 182081 53274 182147 53277
rect 209681 53274 209747 53277
rect 238661 53274 238727 53277
rect 266261 53274 266327 53277
rect 293861 53274 293927 53277
rect 322841 53274 322907 53277
rect 350441 53274 350507 53277
rect 378041 53274 378107 53277
rect 405641 53274 405707 53277
rect 434621 53274 434687 53277
rect 462221 53274 462287 53277
rect 489821 53274 489887 53277
rect 518801 53274 518867 53277
rect 545757 53274 545823 53277
rect 13721 53272 16100 53274
rect 13721 53216 13726 53272
rect 13782 53216 16100 53272
rect 13721 53214 16100 53216
rect 42701 53272 44068 53274
rect 42701 53216 42706 53272
rect 42762 53216 44068 53272
rect 42701 53214 44068 53216
rect 70301 53272 72036 53274
rect 70301 53216 70306 53272
rect 70362 53216 72036 53272
rect 70301 53214 72036 53216
rect 97901 53272 100188 53274
rect 97901 53216 97906 53272
rect 97962 53216 100188 53272
rect 97901 53214 100188 53216
rect 126881 53272 128156 53274
rect 126881 53216 126886 53272
rect 126942 53216 128156 53272
rect 126881 53214 128156 53216
rect 154481 53272 156124 53274
rect 154481 53216 154486 53272
rect 154542 53216 156124 53272
rect 154481 53214 156124 53216
rect 182081 53272 184092 53274
rect 182081 53216 182086 53272
rect 182142 53216 184092 53272
rect 182081 53214 184092 53216
rect 209681 53272 212060 53274
rect 209681 53216 209686 53272
rect 209742 53216 212060 53272
rect 209681 53214 212060 53216
rect 238661 53272 240212 53274
rect 238661 53216 238666 53272
rect 238722 53216 240212 53272
rect 238661 53214 240212 53216
rect 266261 53272 268180 53274
rect 266261 53216 266266 53272
rect 266322 53216 268180 53272
rect 266261 53214 268180 53216
rect 293861 53272 296148 53274
rect 293861 53216 293866 53272
rect 293922 53216 296148 53272
rect 293861 53214 296148 53216
rect 322841 53272 324116 53274
rect 322841 53216 322846 53272
rect 322902 53216 324116 53272
rect 322841 53214 324116 53216
rect 350441 53272 352084 53274
rect 350441 53216 350446 53272
rect 350502 53216 352084 53272
rect 350441 53214 352084 53216
rect 378041 53272 380052 53274
rect 378041 53216 378046 53272
rect 378102 53216 380052 53272
rect 378041 53214 380052 53216
rect 405641 53272 408204 53274
rect 405641 53216 405646 53272
rect 405702 53216 408204 53272
rect 405641 53214 408204 53216
rect 434621 53272 436172 53274
rect 434621 53216 434626 53272
rect 434682 53216 436172 53272
rect 434621 53214 436172 53216
rect 462221 53272 464140 53274
rect 462221 53216 462226 53272
rect 462282 53216 464140 53272
rect 462221 53214 464140 53216
rect 489821 53272 492108 53274
rect 489821 53216 489826 53272
rect 489882 53216 492108 53272
rect 489821 53214 492108 53216
rect 518801 53272 520076 53274
rect 518801 53216 518806 53272
rect 518862 53216 520076 53272
rect 518801 53214 520076 53216
rect 545757 53272 548044 53274
rect 545757 53216 545762 53272
rect 545818 53216 548044 53272
rect 545757 53214 548044 53216
rect 13721 53211 13787 53214
rect 42701 53211 42767 53214
rect 70301 53211 70367 53214
rect 97901 53211 97967 53214
rect 126881 53211 126947 53214
rect 154481 53211 154547 53214
rect 182081 53211 182147 53214
rect 209681 53211 209747 53214
rect 238661 53211 238727 53214
rect 266261 53211 266327 53214
rect 293861 53211 293927 53214
rect 322841 53211 322907 53214
rect 350441 53211 350507 53214
rect 378041 53211 378107 53214
rect 405641 53211 405707 53214
rect 434621 53211 434687 53214
rect 462221 53211 462287 53214
rect 489821 53211 489887 53214
rect 518801 53211 518867 53214
rect 545757 53211 545823 53214
rect 37917 52594 37983 52597
rect 66253 52594 66319 52597
rect 93853 52594 93919 52597
rect 121453 52594 121519 52597
rect 149053 52594 149119 52597
rect 178033 52594 178099 52597
rect 205633 52594 205699 52597
rect 233233 52594 233299 52597
rect 262213 52594 262279 52597
rect 289813 52594 289879 52597
rect 317413 52594 317479 52597
rect 345013 52594 345079 52597
rect 373993 52594 374059 52597
rect 401593 52594 401659 52597
rect 429193 52594 429259 52597
rect 458173 52594 458239 52597
rect 485773 52594 485839 52597
rect 513373 52594 513439 52597
rect 542353 52594 542419 52597
rect 569953 52594 570019 52597
rect 35788 52592 37983 52594
rect 35788 52536 37922 52592
rect 37978 52536 37983 52592
rect 35788 52534 37983 52536
rect 63940 52592 66319 52594
rect 63940 52536 66258 52592
rect 66314 52536 66319 52592
rect 63940 52534 66319 52536
rect 91908 52592 93919 52594
rect 91908 52536 93858 52592
rect 93914 52536 93919 52592
rect 91908 52534 93919 52536
rect 119876 52592 121519 52594
rect 119876 52536 121458 52592
rect 121514 52536 121519 52592
rect 119876 52534 121519 52536
rect 147844 52592 149119 52594
rect 147844 52536 149058 52592
rect 149114 52536 149119 52592
rect 147844 52534 149119 52536
rect 175812 52592 178099 52594
rect 175812 52536 178038 52592
rect 178094 52536 178099 52592
rect 175812 52534 178099 52536
rect 203964 52592 205699 52594
rect 203964 52536 205638 52592
rect 205694 52536 205699 52592
rect 203964 52534 205699 52536
rect 231932 52592 233299 52594
rect 231932 52536 233238 52592
rect 233294 52536 233299 52592
rect 231932 52534 233299 52536
rect 259900 52592 262279 52594
rect 259900 52536 262218 52592
rect 262274 52536 262279 52592
rect 259900 52534 262279 52536
rect 287868 52592 289879 52594
rect 287868 52536 289818 52592
rect 289874 52536 289879 52592
rect 287868 52534 289879 52536
rect 315836 52592 317479 52594
rect 315836 52536 317418 52592
rect 317474 52536 317479 52592
rect 315836 52534 317479 52536
rect 343804 52592 345079 52594
rect 343804 52536 345018 52592
rect 345074 52536 345079 52592
rect 343804 52534 345079 52536
rect 371956 52592 374059 52594
rect 371956 52536 373998 52592
rect 374054 52536 374059 52592
rect 371956 52534 374059 52536
rect 399924 52592 401659 52594
rect 399924 52536 401598 52592
rect 401654 52536 401659 52592
rect 399924 52534 401659 52536
rect 427892 52592 429259 52594
rect 427892 52536 429198 52592
rect 429254 52536 429259 52592
rect 427892 52534 429259 52536
rect 455860 52592 458239 52594
rect 455860 52536 458178 52592
rect 458234 52536 458239 52592
rect 455860 52534 458239 52536
rect 483828 52592 485839 52594
rect 483828 52536 485778 52592
rect 485834 52536 485839 52592
rect 483828 52534 485839 52536
rect 511796 52592 513439 52594
rect 511796 52536 513378 52592
rect 513434 52536 513439 52592
rect 511796 52534 513439 52536
rect 539948 52592 542419 52594
rect 539948 52536 542358 52592
rect 542414 52536 542419 52592
rect 539948 52534 542419 52536
rect 567916 52592 570019 52594
rect 567916 52536 569958 52592
rect 570014 52536 570019 52592
rect 567916 52534 570019 52536
rect 37917 52531 37983 52534
rect 66253 52531 66319 52534
rect 93853 52531 93919 52534
rect 121453 52531 121519 52534
rect 149053 52531 149119 52534
rect 178033 52531 178099 52534
rect 205633 52531 205699 52534
rect 233233 52531 233299 52534
rect 262213 52531 262279 52534
rect 289813 52531 289879 52534
rect 317413 52531 317479 52534
rect 345013 52531 345079 52534
rect 373993 52531 374059 52534
rect 401593 52531 401659 52534
rect 429193 52531 429259 52534
rect 458173 52531 458239 52534
rect 485773 52531 485839 52534
rect 513373 52531 513439 52534
rect 542353 52531 542419 52534
rect 569953 52531 570019 52534
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3233 45522 3299 45525
rect -960 45520 3299 45522
rect -960 45464 3238 45520
rect 3294 45464 3299 45520
rect -960 45462 3299 45464
rect -960 45372 480 45462
rect 3233 45459 3299 45462
rect 61285 36138 61351 36141
rect 61285 36136 61394 36138
rect 61285 36080 61290 36136
rect 61346 36080 61394 36136
rect 61285 36075 61394 36080
rect 11697 35866 11763 35869
rect 11697 35864 16100 35866
rect 11697 35808 11702 35864
rect 11758 35808 16100 35864
rect 61334 35836 61394 36075
rect 11697 35806 16100 35808
rect 11697 35803 11763 35806
rect 63493 33146 63559 33149
rect 61916 33144 63559 33146
rect 61916 33088 63498 33144
rect 63554 33088 63559 33144
rect 61916 33086 63559 33088
rect 63493 33083 63559 33086
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 12433 32466 12499 32469
rect 12433 32464 16100 32466
rect 12433 32408 12438 32464
rect 12494 32408 16100 32464
rect 12433 32406 16100 32408
rect 12433 32403 12499 32406
rect 63585 29746 63651 29749
rect 61916 29744 63651 29746
rect 61916 29688 63590 29744
rect 63646 29688 63651 29744
rect 61916 29686 63651 29688
rect 63585 29683 63651 29686
rect 13721 29066 13787 29069
rect 13721 29064 16100 29066
rect 13721 29008 13726 29064
rect 13782 29008 16100 29064
rect 13721 29006 16100 29008
rect 13721 29003 13787 29006
rect 70301 26890 70367 26893
rect 70301 26888 72066 26890
rect 70301 26832 70306 26888
rect 70362 26832 72066 26888
rect 70301 26830 72066 26832
rect 70301 26827 70367 26830
rect 63493 26346 63559 26349
rect 61916 26344 63559 26346
rect 61916 26288 63498 26344
rect 63554 26288 63559 26344
rect 72006 26316 72066 26830
rect 97901 26346 97967 26349
rect 126881 26346 126947 26349
rect 154481 26346 154547 26349
rect 182081 26346 182147 26349
rect 209681 26346 209747 26349
rect 238661 26346 238727 26349
rect 266261 26346 266327 26349
rect 293861 26346 293927 26349
rect 322841 26346 322907 26349
rect 350441 26346 350507 26349
rect 378041 26346 378107 26349
rect 405641 26346 405707 26349
rect 434621 26346 434687 26349
rect 462221 26346 462287 26349
rect 489821 26346 489887 26349
rect 518801 26346 518867 26349
rect 545757 26346 545823 26349
rect 97901 26344 100188 26346
rect 61916 26286 63559 26288
rect 63493 26283 63559 26286
rect 97901 26288 97906 26344
rect 97962 26288 100188 26344
rect 97901 26286 100188 26288
rect 126881 26344 128156 26346
rect 126881 26288 126886 26344
rect 126942 26288 128156 26344
rect 126881 26286 128156 26288
rect 154481 26344 156124 26346
rect 154481 26288 154486 26344
rect 154542 26288 156124 26344
rect 154481 26286 156124 26288
rect 182081 26344 184092 26346
rect 182081 26288 182086 26344
rect 182142 26288 184092 26344
rect 182081 26286 184092 26288
rect 209681 26344 212060 26346
rect 209681 26288 209686 26344
rect 209742 26288 212060 26344
rect 209681 26286 212060 26288
rect 238661 26344 240212 26346
rect 238661 26288 238666 26344
rect 238722 26288 240212 26344
rect 238661 26286 240212 26288
rect 266261 26344 268180 26346
rect 266261 26288 266266 26344
rect 266322 26288 268180 26344
rect 266261 26286 268180 26288
rect 293861 26344 296148 26346
rect 293861 26288 293866 26344
rect 293922 26288 296148 26344
rect 293861 26286 296148 26288
rect 322841 26344 324116 26346
rect 322841 26288 322846 26344
rect 322902 26288 324116 26344
rect 322841 26286 324116 26288
rect 350441 26344 352084 26346
rect 350441 26288 350446 26344
rect 350502 26288 352084 26344
rect 350441 26286 352084 26288
rect 378041 26344 380052 26346
rect 378041 26288 378046 26344
rect 378102 26288 380052 26344
rect 378041 26286 380052 26288
rect 405641 26344 408204 26346
rect 405641 26288 405646 26344
rect 405702 26288 408204 26344
rect 405641 26286 408204 26288
rect 434621 26344 436172 26346
rect 434621 26288 434626 26344
rect 434682 26288 436172 26344
rect 434621 26286 436172 26288
rect 462221 26344 464140 26346
rect 462221 26288 462226 26344
rect 462282 26288 464140 26344
rect 462221 26286 464140 26288
rect 489821 26344 492108 26346
rect 489821 26288 489826 26344
rect 489882 26288 492108 26344
rect 489821 26286 492108 26288
rect 518801 26344 520076 26346
rect 518801 26288 518806 26344
rect 518862 26288 520076 26344
rect 518801 26286 520076 26288
rect 545757 26344 548044 26346
rect 545757 26288 545762 26344
rect 545818 26288 548044 26344
rect 545757 26286 548044 26288
rect 97901 26283 97967 26286
rect 126881 26283 126947 26286
rect 154481 26283 154547 26286
rect 182081 26283 182147 26286
rect 209681 26283 209747 26286
rect 238661 26283 238727 26286
rect 266261 26283 266327 26286
rect 293861 26283 293927 26286
rect 322841 26283 322907 26286
rect 350441 26283 350507 26286
rect 378041 26283 378107 26286
rect 405641 26283 405707 26286
rect 434621 26283 434687 26286
rect 462221 26283 462287 26286
rect 489821 26283 489887 26286
rect 518801 26283 518867 26286
rect 545757 26283 545823 26286
rect 205633 25938 205699 25941
rect 203934 25936 205699 25938
rect 203934 25880 205638 25936
rect 205694 25880 205699 25936
rect 203934 25878 205699 25880
rect 13721 25666 13787 25669
rect 93853 25666 93919 25669
rect 121453 25666 121519 25669
rect 149053 25666 149119 25669
rect 178033 25666 178099 25669
rect 13721 25664 16100 25666
rect 13721 25608 13726 25664
rect 13782 25608 16100 25664
rect 13721 25606 16100 25608
rect 91908 25664 93919 25666
rect 91908 25608 93858 25664
rect 93914 25608 93919 25664
rect 91908 25606 93919 25608
rect 119876 25664 121519 25666
rect 119876 25608 121458 25664
rect 121514 25608 121519 25664
rect 119876 25606 121519 25608
rect 147844 25664 149119 25666
rect 147844 25608 149058 25664
rect 149114 25608 149119 25664
rect 147844 25606 149119 25608
rect 175812 25664 178099 25666
rect 175812 25608 178038 25664
rect 178094 25608 178099 25664
rect 203934 25636 203994 25878
rect 205633 25875 205699 25878
rect 233233 25666 233299 25669
rect 262213 25666 262279 25669
rect 289813 25666 289879 25669
rect 317413 25666 317479 25669
rect 345013 25666 345079 25669
rect 373993 25666 374059 25669
rect 401593 25666 401659 25669
rect 429193 25666 429259 25669
rect 458173 25666 458239 25669
rect 485773 25666 485839 25669
rect 513373 25666 513439 25669
rect 542353 25666 542419 25669
rect 569953 25666 570019 25669
rect 231932 25664 233299 25666
rect 175812 25606 178099 25608
rect 231932 25608 233238 25664
rect 233294 25608 233299 25664
rect 231932 25606 233299 25608
rect 259900 25664 262279 25666
rect 259900 25608 262218 25664
rect 262274 25608 262279 25664
rect 259900 25606 262279 25608
rect 287868 25664 289879 25666
rect 287868 25608 289818 25664
rect 289874 25608 289879 25664
rect 287868 25606 289879 25608
rect 315836 25664 317479 25666
rect 315836 25608 317418 25664
rect 317474 25608 317479 25664
rect 315836 25606 317479 25608
rect 343804 25664 345079 25666
rect 343804 25608 345018 25664
rect 345074 25608 345079 25664
rect 343804 25606 345079 25608
rect 371956 25664 374059 25666
rect 371956 25608 373998 25664
rect 374054 25608 374059 25664
rect 371956 25606 374059 25608
rect 399924 25664 401659 25666
rect 399924 25608 401598 25664
rect 401654 25608 401659 25664
rect 399924 25606 401659 25608
rect 427892 25664 429259 25666
rect 427892 25608 429198 25664
rect 429254 25608 429259 25664
rect 427892 25606 429259 25608
rect 455860 25664 458239 25666
rect 455860 25608 458178 25664
rect 458234 25608 458239 25664
rect 455860 25606 458239 25608
rect 483828 25664 485839 25666
rect 483828 25608 485778 25664
rect 485834 25608 485839 25664
rect 483828 25606 485839 25608
rect 511796 25664 513439 25666
rect 511796 25608 513378 25664
rect 513434 25608 513439 25664
rect 511796 25606 513439 25608
rect 539948 25664 542419 25666
rect 539948 25608 542358 25664
rect 542414 25608 542419 25664
rect 539948 25606 542419 25608
rect 567916 25664 570019 25666
rect 567916 25608 569958 25664
rect 570014 25608 570019 25664
rect 567916 25606 570019 25608
rect 13721 25603 13787 25606
rect 93853 25603 93919 25606
rect 121453 25603 121519 25606
rect 149053 25603 149119 25606
rect 178033 25603 178099 25606
rect 233233 25603 233299 25606
rect 262213 25603 262279 25606
rect 289813 25603 289879 25606
rect 317413 25603 317479 25606
rect 345013 25603 345079 25606
rect 373993 25603 374059 25606
rect 401593 25603 401659 25606
rect 429193 25603 429259 25606
rect 458173 25603 458239 25606
rect 485773 25603 485839 25606
rect 513373 25603 513439 25606
rect 542353 25603 542419 25606
rect 569953 25603 570019 25606
rect 64229 22946 64295 22949
rect 61916 22944 64295 22946
rect 61916 22888 64234 22944
rect 64290 22888 64295 22944
rect 61916 22886 64295 22888
rect 64229 22883 64295 22886
rect 13169 22266 13235 22269
rect 13169 22264 16100 22266
rect 13169 22208 13174 22264
rect 13230 22208 16100 22264
rect 13169 22206 16100 22208
rect 13169 22203 13235 22206
rect 583520 19668 584960 19908
rect 63493 19546 63559 19549
rect 61916 19544 63559 19546
rect -960 19410 480 19500
rect 61916 19488 63498 19544
rect 63554 19488 63559 19544
rect 61916 19486 63559 19488
rect 63493 19483 63559 19486
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 12433 18866 12499 18869
rect 12433 18864 16100 18866
rect 12433 18808 12438 18864
rect 12494 18808 16100 18864
rect 12433 18806 16100 18808
rect 12433 18803 12499 18806
rect 64413 16146 64479 16149
rect 61916 16144 64479 16146
rect 61916 16088 64418 16144
rect 64474 16088 64479 16144
rect 61916 16086 64479 16088
rect 64413 16083 64479 16086
rect -960 6490 480 6580
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6716
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 698454 -2346 705242
rect 37994 705798 38614 711590
rect 37994 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 38614 705798
rect 37994 705478 38614 705562
rect 37994 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 38614 705478
rect -2966 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 -2346 698454
rect -2966 698134 -2346 698218
rect -2966 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 -2346 698134
rect -2966 671454 -2346 697898
rect -2966 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 -2346 671454
rect -2966 671134 -2346 671218
rect -2966 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 -2346 671134
rect -2966 644454 -2346 670898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 617454 -2346 643898
rect -2966 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 -2346 617454
rect -2966 617134 -2346 617218
rect -2966 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 -2346 617134
rect -2966 590454 -2346 616898
rect -2966 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 -2346 590454
rect -2966 590134 -2346 590218
rect -2966 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 -2346 590134
rect -2966 563454 -2346 589898
rect -2966 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 -2346 563454
rect -2966 563134 -2346 563218
rect -2966 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 -2346 563134
rect -2966 536454 -2346 562898
rect -2966 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 -2346 536454
rect -2966 536134 -2346 536218
rect -2966 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 -2346 536134
rect -2966 509454 -2346 535898
rect -2966 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 -2346 509454
rect -2966 509134 -2346 509218
rect -2966 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 -2346 509134
rect -2966 482454 -2346 508898
rect -2966 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 -2346 482454
rect -2966 482134 -2346 482218
rect -2966 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 -2346 482134
rect -2966 455454 -2346 481898
rect -2966 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 -2346 455454
rect -2966 455134 -2346 455218
rect -2966 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 -2346 455134
rect -2966 428454 -2346 454898
rect -2966 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 -2346 428454
rect -2966 428134 -2346 428218
rect -2966 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 -2346 428134
rect -2966 401454 -2346 427898
rect -2966 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 -2346 401454
rect -2966 401134 -2346 401218
rect -2966 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 -2346 401134
rect -2966 374454 -2346 400898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 347454 -2346 373898
rect -2966 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 -2346 347454
rect -2966 347134 -2346 347218
rect -2966 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 -2346 347134
rect -2966 320454 -2346 346898
rect -2966 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 -2346 320454
rect -2966 320134 -2346 320218
rect -2966 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 -2346 320134
rect -2966 293454 -2346 319898
rect -2966 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 -2346 293454
rect -2966 293134 -2346 293218
rect -2966 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 -2346 293134
rect -2966 266454 -2346 292898
rect -2966 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 -2346 266454
rect -2966 266134 -2346 266218
rect -2966 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 -2346 266134
rect -2966 239454 -2346 265898
rect -2966 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 -2346 239454
rect -2966 239134 -2346 239218
rect -2966 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 -2346 239134
rect -2966 212454 -2346 238898
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 -2346 212454
rect -2966 212134 -2346 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 -2346 212134
rect -2966 185454 -2346 211898
rect -2966 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 -2346 185454
rect -2966 185134 -2346 185218
rect -2966 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 -2346 185134
rect -2966 158454 -2346 184898
rect -2966 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 -2346 158454
rect -2966 158134 -2346 158218
rect -2966 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 -2346 158134
rect -2966 131454 -2346 157898
rect -2966 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 -2346 131454
rect -2966 131134 -2346 131218
rect -2966 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 -2346 131134
rect -2966 104454 -2346 130898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 77454 -2346 103898
rect -2966 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 -2346 77454
rect -2966 77134 -2346 77218
rect -2966 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 -2346 77134
rect -2966 50454 -2346 76898
rect -2966 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 -2346 50454
rect -2966 50134 -2346 50218
rect -2966 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 -2346 50134
rect -2966 23454 -2346 49898
rect -2966 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 -2346 23454
rect -2966 23134 -2346 23218
rect -2966 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 -2346 23134
rect -2966 -1306 -2346 22898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 701829 -1386 704282
rect -2006 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 -1386 701829
rect -2006 701509 -1386 701593
rect -2006 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 -1386 701509
rect -2006 674829 -1386 701273
rect 37994 698454 38614 705242
rect 37994 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 38614 698454
rect 37994 698134 38614 698218
rect 37994 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 38614 698134
rect 37994 686000 38614 697898
rect 41494 704838 42114 711590
rect 41494 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 42114 704838
rect 41494 704518 42114 704602
rect 41494 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 42114 704518
rect 41494 701829 42114 704282
rect 41494 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 42114 701829
rect 41494 701509 42114 701593
rect 41494 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 42114 701509
rect 41494 686000 42114 701273
rect 65994 705798 66614 711590
rect 65994 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 66614 705798
rect 65994 705478 66614 705562
rect 65994 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 66614 705478
rect 65994 698454 66614 705242
rect 65994 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 66614 698454
rect 65994 698134 66614 698218
rect 65994 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 66614 698134
rect 65994 686000 66614 697898
rect 69494 704838 70114 711590
rect 69494 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 70114 704838
rect 69494 704518 70114 704602
rect 69494 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 70114 704518
rect 69494 701829 70114 704282
rect 69494 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 70114 701829
rect 69494 701509 70114 701593
rect 69494 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 70114 701509
rect 69494 686000 70114 701273
rect 93994 705798 94614 711590
rect 93994 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 94614 705798
rect 93994 705478 94614 705562
rect 93994 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 94614 705478
rect 93994 698454 94614 705242
rect 93994 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 94614 698454
rect 93994 698134 94614 698218
rect 93994 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 94614 698134
rect 93994 686000 94614 697898
rect 97494 704838 98114 711590
rect 97494 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 98114 704838
rect 97494 704518 98114 704602
rect 97494 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 98114 704518
rect 97494 701829 98114 704282
rect 97494 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 98114 701829
rect 97494 701509 98114 701593
rect 97494 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 98114 701509
rect 97494 686000 98114 701273
rect 121994 705798 122614 711590
rect 121994 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 122614 705798
rect 121994 705478 122614 705562
rect 121994 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 122614 705478
rect 121994 698454 122614 705242
rect 121994 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 122614 698454
rect 121994 698134 122614 698218
rect 121994 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 122614 698134
rect 121994 686000 122614 697898
rect 125494 704838 126114 711590
rect 125494 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 126114 704838
rect 125494 704518 126114 704602
rect 125494 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 126114 704518
rect 125494 701829 126114 704282
rect 125494 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 126114 701829
rect 125494 701509 126114 701593
rect 125494 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 126114 701509
rect 125494 686000 126114 701273
rect 149994 705798 150614 711590
rect 149994 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 150614 705798
rect 149994 705478 150614 705562
rect 149994 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 150614 705478
rect 149994 698454 150614 705242
rect 149994 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 150614 698454
rect 149994 698134 150614 698218
rect 149994 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 150614 698134
rect 149994 686000 150614 697898
rect 153494 704838 154114 711590
rect 153494 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 154114 704838
rect 153494 704518 154114 704602
rect 153494 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 154114 704518
rect 153494 701829 154114 704282
rect 153494 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 154114 701829
rect 153494 701509 154114 701593
rect 153494 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 154114 701509
rect 153494 686000 154114 701273
rect 177994 705798 178614 711590
rect 177994 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 178614 705798
rect 177994 705478 178614 705562
rect 177994 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 178614 705478
rect 177994 698454 178614 705242
rect 177994 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 178614 698454
rect 177994 698134 178614 698218
rect 177994 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 178614 698134
rect 177994 686000 178614 697898
rect 181494 704838 182114 711590
rect 181494 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 182114 704838
rect 181494 704518 182114 704602
rect 181494 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 182114 704518
rect 181494 701829 182114 704282
rect 181494 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 182114 701829
rect 181494 701509 182114 701593
rect 181494 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 182114 701509
rect 181494 686000 182114 701273
rect 205994 705798 206614 711590
rect 205994 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 206614 705798
rect 205994 705478 206614 705562
rect 205994 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 206614 705478
rect 205994 698454 206614 705242
rect 205994 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 206614 698454
rect 205994 698134 206614 698218
rect 205994 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 206614 698134
rect 205994 686000 206614 697898
rect 209494 704838 210114 711590
rect 209494 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 210114 704838
rect 209494 704518 210114 704602
rect 209494 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 210114 704518
rect 209494 701829 210114 704282
rect 209494 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 210114 701829
rect 209494 701509 210114 701593
rect 209494 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 210114 701509
rect 209494 686000 210114 701273
rect 233994 705798 234614 711590
rect 233994 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 234614 705798
rect 233994 705478 234614 705562
rect 233994 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 234614 705478
rect 233994 698454 234614 705242
rect 233994 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 234614 698454
rect 233994 698134 234614 698218
rect 233994 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 234614 698134
rect 233994 686000 234614 697898
rect 237494 704838 238114 711590
rect 237494 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 238114 704838
rect 237494 704518 238114 704602
rect 237494 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 238114 704518
rect 237494 701829 238114 704282
rect 237494 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 238114 701829
rect 237494 701509 238114 701593
rect 237494 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 238114 701509
rect 237494 686000 238114 701273
rect 261994 705798 262614 711590
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 698454 262614 705242
rect 261994 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 262614 698454
rect 261994 698134 262614 698218
rect 261994 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 262614 698134
rect 261994 686000 262614 697898
rect 265494 704838 266114 711590
rect 265494 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 266114 704838
rect 265494 704518 266114 704602
rect 265494 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 266114 704518
rect 265494 701829 266114 704282
rect 265494 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 266114 701829
rect 265494 701509 266114 701593
rect 265494 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 266114 701509
rect 265494 686000 266114 701273
rect 289994 705798 290614 711590
rect 289994 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 290614 705798
rect 289994 705478 290614 705562
rect 289994 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 290614 705478
rect 289994 698454 290614 705242
rect 289994 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 290614 698454
rect 289994 698134 290614 698218
rect 289994 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 290614 698134
rect 289994 686000 290614 697898
rect 293494 704838 294114 711590
rect 293494 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 294114 704838
rect 293494 704518 294114 704602
rect 293494 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 294114 704518
rect 293494 701829 294114 704282
rect 293494 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 294114 701829
rect 293494 701509 294114 701593
rect 293494 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 294114 701509
rect 293494 686000 294114 701273
rect 317994 705798 318614 711590
rect 317994 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 318614 705798
rect 317994 705478 318614 705562
rect 317994 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 318614 705478
rect 317994 698454 318614 705242
rect 317994 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 318614 698454
rect 317994 698134 318614 698218
rect 317994 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 318614 698134
rect 317994 686000 318614 697898
rect 321494 704838 322114 711590
rect 321494 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 322114 704838
rect 321494 704518 322114 704602
rect 321494 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 322114 704518
rect 321494 701829 322114 704282
rect 321494 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 322114 701829
rect 321494 701509 322114 701593
rect 321494 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 322114 701509
rect 321494 686000 322114 701273
rect 345994 705798 346614 711590
rect 345994 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 346614 705798
rect 345994 705478 346614 705562
rect 345994 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 346614 705478
rect 345994 698454 346614 705242
rect 345994 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 346614 698454
rect 345994 698134 346614 698218
rect 345994 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 346614 698134
rect 345994 686000 346614 697898
rect 349494 704838 350114 711590
rect 349494 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 350114 704838
rect 349494 704518 350114 704602
rect 349494 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 350114 704518
rect 349494 701829 350114 704282
rect 349494 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 350114 701829
rect 349494 701509 350114 701593
rect 349494 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 350114 701509
rect 349494 686000 350114 701273
rect 373994 705798 374614 711590
rect 373994 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 374614 705798
rect 373994 705478 374614 705562
rect 373994 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 374614 705478
rect 373994 698454 374614 705242
rect 373994 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 374614 698454
rect 373994 698134 374614 698218
rect 373994 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 374614 698134
rect 373994 686000 374614 697898
rect 377494 704838 378114 711590
rect 377494 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 378114 704838
rect 377494 704518 378114 704602
rect 377494 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 378114 704518
rect 377494 701829 378114 704282
rect 377494 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 378114 701829
rect 377494 701509 378114 701593
rect 377494 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 378114 701509
rect 377494 686000 378114 701273
rect 401994 705798 402614 711590
rect 401994 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 402614 705798
rect 401994 705478 402614 705562
rect 401994 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 402614 705478
rect 401994 698454 402614 705242
rect 401994 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 402614 698454
rect 401994 698134 402614 698218
rect 401994 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 402614 698134
rect 401994 686000 402614 697898
rect 405494 704838 406114 711590
rect 405494 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 406114 704838
rect 405494 704518 406114 704602
rect 405494 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 406114 704518
rect 405494 701829 406114 704282
rect 405494 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 406114 701829
rect 405494 701509 406114 701593
rect 405494 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 406114 701509
rect 405494 686000 406114 701273
rect 429994 705798 430614 711590
rect 429994 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 430614 705798
rect 429994 705478 430614 705562
rect 429994 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 430614 705478
rect 429994 698454 430614 705242
rect 429994 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 430614 698454
rect 429994 698134 430614 698218
rect 429994 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 430614 698134
rect 429994 686000 430614 697898
rect 433494 704838 434114 711590
rect 433494 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 434114 704838
rect 433494 704518 434114 704602
rect 433494 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 434114 704518
rect 433494 701829 434114 704282
rect 433494 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 434114 701829
rect 433494 701509 434114 701593
rect 433494 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 434114 701509
rect 433494 686000 434114 701273
rect 457994 705798 458614 711590
rect 457994 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 458614 705798
rect 457994 705478 458614 705562
rect 457994 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 458614 705478
rect 457994 698454 458614 705242
rect 457994 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 458614 698454
rect 457994 698134 458614 698218
rect 457994 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 458614 698134
rect 457994 686000 458614 697898
rect 461494 704838 462114 711590
rect 461494 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 462114 704838
rect 461494 704518 462114 704602
rect 461494 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 462114 704518
rect 461494 701829 462114 704282
rect 461494 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 462114 701829
rect 461494 701509 462114 701593
rect 461494 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 462114 701509
rect 461494 686000 462114 701273
rect 485994 705798 486614 711590
rect 485994 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 486614 705798
rect 485994 705478 486614 705562
rect 485994 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 486614 705478
rect 485994 698454 486614 705242
rect 485994 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 486614 698454
rect 485994 698134 486614 698218
rect 485994 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 486614 698134
rect 485994 686000 486614 697898
rect 489494 704838 490114 711590
rect 489494 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 490114 704838
rect 489494 704518 490114 704602
rect 489494 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 490114 704518
rect 489494 701829 490114 704282
rect 489494 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 490114 701829
rect 489494 701509 490114 701593
rect 489494 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 490114 701509
rect 489494 686000 490114 701273
rect 513994 705798 514614 711590
rect 513994 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 514614 705798
rect 513994 705478 514614 705562
rect 513994 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 514614 705478
rect 513994 698454 514614 705242
rect 513994 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 514614 698454
rect 513994 698134 514614 698218
rect 513994 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 514614 698134
rect 513994 686000 514614 697898
rect 517494 704838 518114 711590
rect 517494 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 518114 704838
rect 517494 704518 518114 704602
rect 517494 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 518114 704518
rect 517494 701829 518114 704282
rect 517494 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 518114 701829
rect 517494 701509 518114 701593
rect 517494 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 518114 701509
rect 517494 686000 518114 701273
rect 541994 705798 542614 711590
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 541994 698454 542614 705242
rect 541994 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 542614 698454
rect 541994 698134 542614 698218
rect 541994 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 542614 698134
rect 541994 686000 542614 697898
rect 545494 704838 546114 711590
rect 545494 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 546114 704838
rect 545494 704518 546114 704602
rect 545494 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 546114 704518
rect 545494 701829 546114 704282
rect 545494 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 546114 701829
rect 545494 701509 546114 701593
rect 545494 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 546114 701509
rect 545494 686000 546114 701273
rect 569994 705798 570614 711590
rect 569994 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 570614 705798
rect 569994 705478 570614 705562
rect 569994 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 570614 705478
rect 569994 698454 570614 705242
rect 569994 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 570614 698454
rect 569994 698134 570614 698218
rect 569994 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 570614 698134
rect 569994 686000 570614 697898
rect 573494 704838 574114 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 573494 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 574114 704838
rect 573494 704518 574114 704602
rect 573494 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 574114 704518
rect 573494 701829 574114 704282
rect 573494 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 574114 701829
rect 573494 701509 574114 701593
rect 573494 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 574114 701509
rect -2006 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 -1386 674829
rect -2006 674509 -1386 674593
rect -2006 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 -1386 674509
rect -2006 647829 -1386 674273
rect 19910 674829 20230 674861
rect 19910 674593 19952 674829
rect 20188 674593 20230 674829
rect 19910 674509 20230 674593
rect 19910 674273 19952 674509
rect 20188 674273 20230 674509
rect 19910 674241 20230 674273
rect 25840 674829 26160 674861
rect 25840 674593 25882 674829
rect 26118 674593 26160 674829
rect 25840 674509 26160 674593
rect 25840 674273 25882 674509
rect 26118 674273 26160 674509
rect 25840 674241 26160 674273
rect 31771 674829 32091 674861
rect 31771 674593 31813 674829
rect 32049 674593 32091 674829
rect 31771 674509 32091 674593
rect 31771 674273 31813 674509
rect 32049 674273 32091 674509
rect 31771 674241 32091 674273
rect 47910 674829 48230 674861
rect 47910 674593 47952 674829
rect 48188 674593 48230 674829
rect 47910 674509 48230 674593
rect 47910 674273 47952 674509
rect 48188 674273 48230 674509
rect 47910 674241 48230 674273
rect 53840 674829 54160 674861
rect 53840 674593 53882 674829
rect 54118 674593 54160 674829
rect 53840 674509 54160 674593
rect 53840 674273 53882 674509
rect 54118 674273 54160 674509
rect 53840 674241 54160 674273
rect 59771 674829 60091 674861
rect 59771 674593 59813 674829
rect 60049 674593 60091 674829
rect 59771 674509 60091 674593
rect 59771 674273 59813 674509
rect 60049 674273 60091 674509
rect 59771 674241 60091 674273
rect 75910 674829 76230 674861
rect 75910 674593 75952 674829
rect 76188 674593 76230 674829
rect 75910 674509 76230 674593
rect 75910 674273 75952 674509
rect 76188 674273 76230 674509
rect 75910 674241 76230 674273
rect 81840 674829 82160 674861
rect 81840 674593 81882 674829
rect 82118 674593 82160 674829
rect 81840 674509 82160 674593
rect 81840 674273 81882 674509
rect 82118 674273 82160 674509
rect 81840 674241 82160 674273
rect 87771 674829 88091 674861
rect 87771 674593 87813 674829
rect 88049 674593 88091 674829
rect 87771 674509 88091 674593
rect 87771 674273 87813 674509
rect 88049 674273 88091 674509
rect 87771 674241 88091 674273
rect 103910 674829 104230 674861
rect 103910 674593 103952 674829
rect 104188 674593 104230 674829
rect 103910 674509 104230 674593
rect 103910 674273 103952 674509
rect 104188 674273 104230 674509
rect 103910 674241 104230 674273
rect 109840 674829 110160 674861
rect 109840 674593 109882 674829
rect 110118 674593 110160 674829
rect 109840 674509 110160 674593
rect 109840 674273 109882 674509
rect 110118 674273 110160 674509
rect 109840 674241 110160 674273
rect 115771 674829 116091 674861
rect 115771 674593 115813 674829
rect 116049 674593 116091 674829
rect 115771 674509 116091 674593
rect 115771 674273 115813 674509
rect 116049 674273 116091 674509
rect 115771 674241 116091 674273
rect 131910 674829 132230 674861
rect 131910 674593 131952 674829
rect 132188 674593 132230 674829
rect 131910 674509 132230 674593
rect 131910 674273 131952 674509
rect 132188 674273 132230 674509
rect 131910 674241 132230 674273
rect 137840 674829 138160 674861
rect 137840 674593 137882 674829
rect 138118 674593 138160 674829
rect 137840 674509 138160 674593
rect 137840 674273 137882 674509
rect 138118 674273 138160 674509
rect 137840 674241 138160 674273
rect 143771 674829 144091 674861
rect 143771 674593 143813 674829
rect 144049 674593 144091 674829
rect 143771 674509 144091 674593
rect 143771 674273 143813 674509
rect 144049 674273 144091 674509
rect 143771 674241 144091 674273
rect 159910 674829 160230 674861
rect 159910 674593 159952 674829
rect 160188 674593 160230 674829
rect 159910 674509 160230 674593
rect 159910 674273 159952 674509
rect 160188 674273 160230 674509
rect 159910 674241 160230 674273
rect 165840 674829 166160 674861
rect 165840 674593 165882 674829
rect 166118 674593 166160 674829
rect 165840 674509 166160 674593
rect 165840 674273 165882 674509
rect 166118 674273 166160 674509
rect 165840 674241 166160 674273
rect 171771 674829 172091 674861
rect 171771 674593 171813 674829
rect 172049 674593 172091 674829
rect 171771 674509 172091 674593
rect 171771 674273 171813 674509
rect 172049 674273 172091 674509
rect 171771 674241 172091 674273
rect 187910 674829 188230 674861
rect 187910 674593 187952 674829
rect 188188 674593 188230 674829
rect 187910 674509 188230 674593
rect 187910 674273 187952 674509
rect 188188 674273 188230 674509
rect 187910 674241 188230 674273
rect 193840 674829 194160 674861
rect 193840 674593 193882 674829
rect 194118 674593 194160 674829
rect 193840 674509 194160 674593
rect 193840 674273 193882 674509
rect 194118 674273 194160 674509
rect 193840 674241 194160 674273
rect 199771 674829 200091 674861
rect 199771 674593 199813 674829
rect 200049 674593 200091 674829
rect 199771 674509 200091 674593
rect 199771 674273 199813 674509
rect 200049 674273 200091 674509
rect 199771 674241 200091 674273
rect 215910 674829 216230 674861
rect 215910 674593 215952 674829
rect 216188 674593 216230 674829
rect 215910 674509 216230 674593
rect 215910 674273 215952 674509
rect 216188 674273 216230 674509
rect 215910 674241 216230 674273
rect 221840 674829 222160 674861
rect 221840 674593 221882 674829
rect 222118 674593 222160 674829
rect 221840 674509 222160 674593
rect 221840 674273 221882 674509
rect 222118 674273 222160 674509
rect 221840 674241 222160 674273
rect 227771 674829 228091 674861
rect 227771 674593 227813 674829
rect 228049 674593 228091 674829
rect 227771 674509 228091 674593
rect 227771 674273 227813 674509
rect 228049 674273 228091 674509
rect 227771 674241 228091 674273
rect 243910 674829 244230 674861
rect 243910 674593 243952 674829
rect 244188 674593 244230 674829
rect 243910 674509 244230 674593
rect 243910 674273 243952 674509
rect 244188 674273 244230 674509
rect 243910 674241 244230 674273
rect 249840 674829 250160 674861
rect 249840 674593 249882 674829
rect 250118 674593 250160 674829
rect 249840 674509 250160 674593
rect 249840 674273 249882 674509
rect 250118 674273 250160 674509
rect 249840 674241 250160 674273
rect 255771 674829 256091 674861
rect 255771 674593 255813 674829
rect 256049 674593 256091 674829
rect 255771 674509 256091 674593
rect 255771 674273 255813 674509
rect 256049 674273 256091 674509
rect 255771 674241 256091 674273
rect 271910 674829 272230 674861
rect 271910 674593 271952 674829
rect 272188 674593 272230 674829
rect 271910 674509 272230 674593
rect 271910 674273 271952 674509
rect 272188 674273 272230 674509
rect 271910 674241 272230 674273
rect 277840 674829 278160 674861
rect 277840 674593 277882 674829
rect 278118 674593 278160 674829
rect 277840 674509 278160 674593
rect 277840 674273 277882 674509
rect 278118 674273 278160 674509
rect 277840 674241 278160 674273
rect 283771 674829 284091 674861
rect 283771 674593 283813 674829
rect 284049 674593 284091 674829
rect 283771 674509 284091 674593
rect 283771 674273 283813 674509
rect 284049 674273 284091 674509
rect 283771 674241 284091 674273
rect 299910 674829 300230 674861
rect 299910 674593 299952 674829
rect 300188 674593 300230 674829
rect 299910 674509 300230 674593
rect 299910 674273 299952 674509
rect 300188 674273 300230 674509
rect 299910 674241 300230 674273
rect 305840 674829 306160 674861
rect 305840 674593 305882 674829
rect 306118 674593 306160 674829
rect 305840 674509 306160 674593
rect 305840 674273 305882 674509
rect 306118 674273 306160 674509
rect 305840 674241 306160 674273
rect 311771 674829 312091 674861
rect 311771 674593 311813 674829
rect 312049 674593 312091 674829
rect 311771 674509 312091 674593
rect 311771 674273 311813 674509
rect 312049 674273 312091 674509
rect 311771 674241 312091 674273
rect 327910 674829 328230 674861
rect 327910 674593 327952 674829
rect 328188 674593 328230 674829
rect 327910 674509 328230 674593
rect 327910 674273 327952 674509
rect 328188 674273 328230 674509
rect 327910 674241 328230 674273
rect 333840 674829 334160 674861
rect 333840 674593 333882 674829
rect 334118 674593 334160 674829
rect 333840 674509 334160 674593
rect 333840 674273 333882 674509
rect 334118 674273 334160 674509
rect 333840 674241 334160 674273
rect 339771 674829 340091 674861
rect 339771 674593 339813 674829
rect 340049 674593 340091 674829
rect 339771 674509 340091 674593
rect 339771 674273 339813 674509
rect 340049 674273 340091 674509
rect 339771 674241 340091 674273
rect 355910 674829 356230 674861
rect 355910 674593 355952 674829
rect 356188 674593 356230 674829
rect 355910 674509 356230 674593
rect 355910 674273 355952 674509
rect 356188 674273 356230 674509
rect 355910 674241 356230 674273
rect 361840 674829 362160 674861
rect 361840 674593 361882 674829
rect 362118 674593 362160 674829
rect 361840 674509 362160 674593
rect 361840 674273 361882 674509
rect 362118 674273 362160 674509
rect 361840 674241 362160 674273
rect 367771 674829 368091 674861
rect 367771 674593 367813 674829
rect 368049 674593 368091 674829
rect 367771 674509 368091 674593
rect 367771 674273 367813 674509
rect 368049 674273 368091 674509
rect 367771 674241 368091 674273
rect 383910 674829 384230 674861
rect 383910 674593 383952 674829
rect 384188 674593 384230 674829
rect 383910 674509 384230 674593
rect 383910 674273 383952 674509
rect 384188 674273 384230 674509
rect 383910 674241 384230 674273
rect 389840 674829 390160 674861
rect 389840 674593 389882 674829
rect 390118 674593 390160 674829
rect 389840 674509 390160 674593
rect 389840 674273 389882 674509
rect 390118 674273 390160 674509
rect 389840 674241 390160 674273
rect 395771 674829 396091 674861
rect 395771 674593 395813 674829
rect 396049 674593 396091 674829
rect 395771 674509 396091 674593
rect 395771 674273 395813 674509
rect 396049 674273 396091 674509
rect 395771 674241 396091 674273
rect 411910 674829 412230 674861
rect 411910 674593 411952 674829
rect 412188 674593 412230 674829
rect 411910 674509 412230 674593
rect 411910 674273 411952 674509
rect 412188 674273 412230 674509
rect 411910 674241 412230 674273
rect 417840 674829 418160 674861
rect 417840 674593 417882 674829
rect 418118 674593 418160 674829
rect 417840 674509 418160 674593
rect 417840 674273 417882 674509
rect 418118 674273 418160 674509
rect 417840 674241 418160 674273
rect 423771 674829 424091 674861
rect 423771 674593 423813 674829
rect 424049 674593 424091 674829
rect 423771 674509 424091 674593
rect 423771 674273 423813 674509
rect 424049 674273 424091 674509
rect 423771 674241 424091 674273
rect 439910 674829 440230 674861
rect 439910 674593 439952 674829
rect 440188 674593 440230 674829
rect 439910 674509 440230 674593
rect 439910 674273 439952 674509
rect 440188 674273 440230 674509
rect 439910 674241 440230 674273
rect 445840 674829 446160 674861
rect 445840 674593 445882 674829
rect 446118 674593 446160 674829
rect 445840 674509 446160 674593
rect 445840 674273 445882 674509
rect 446118 674273 446160 674509
rect 445840 674241 446160 674273
rect 451771 674829 452091 674861
rect 451771 674593 451813 674829
rect 452049 674593 452091 674829
rect 451771 674509 452091 674593
rect 451771 674273 451813 674509
rect 452049 674273 452091 674509
rect 451771 674241 452091 674273
rect 467910 674829 468230 674861
rect 467910 674593 467952 674829
rect 468188 674593 468230 674829
rect 467910 674509 468230 674593
rect 467910 674273 467952 674509
rect 468188 674273 468230 674509
rect 467910 674241 468230 674273
rect 473840 674829 474160 674861
rect 473840 674593 473882 674829
rect 474118 674593 474160 674829
rect 473840 674509 474160 674593
rect 473840 674273 473882 674509
rect 474118 674273 474160 674509
rect 473840 674241 474160 674273
rect 479771 674829 480091 674861
rect 479771 674593 479813 674829
rect 480049 674593 480091 674829
rect 479771 674509 480091 674593
rect 479771 674273 479813 674509
rect 480049 674273 480091 674509
rect 479771 674241 480091 674273
rect 495910 674829 496230 674861
rect 495910 674593 495952 674829
rect 496188 674593 496230 674829
rect 495910 674509 496230 674593
rect 495910 674273 495952 674509
rect 496188 674273 496230 674509
rect 495910 674241 496230 674273
rect 501840 674829 502160 674861
rect 501840 674593 501882 674829
rect 502118 674593 502160 674829
rect 501840 674509 502160 674593
rect 501840 674273 501882 674509
rect 502118 674273 502160 674509
rect 501840 674241 502160 674273
rect 507771 674829 508091 674861
rect 507771 674593 507813 674829
rect 508049 674593 508091 674829
rect 507771 674509 508091 674593
rect 507771 674273 507813 674509
rect 508049 674273 508091 674509
rect 507771 674241 508091 674273
rect 523910 674829 524230 674861
rect 523910 674593 523952 674829
rect 524188 674593 524230 674829
rect 523910 674509 524230 674593
rect 523910 674273 523952 674509
rect 524188 674273 524230 674509
rect 523910 674241 524230 674273
rect 529840 674829 530160 674861
rect 529840 674593 529882 674829
rect 530118 674593 530160 674829
rect 529840 674509 530160 674593
rect 529840 674273 529882 674509
rect 530118 674273 530160 674509
rect 529840 674241 530160 674273
rect 535771 674829 536091 674861
rect 535771 674593 535813 674829
rect 536049 674593 536091 674829
rect 535771 674509 536091 674593
rect 535771 674273 535813 674509
rect 536049 674273 536091 674509
rect 535771 674241 536091 674273
rect 551910 674829 552230 674861
rect 551910 674593 551952 674829
rect 552188 674593 552230 674829
rect 551910 674509 552230 674593
rect 551910 674273 551952 674509
rect 552188 674273 552230 674509
rect 551910 674241 552230 674273
rect 557840 674829 558160 674861
rect 557840 674593 557882 674829
rect 558118 674593 558160 674829
rect 557840 674509 558160 674593
rect 557840 674273 557882 674509
rect 558118 674273 558160 674509
rect 557840 674241 558160 674273
rect 563771 674829 564091 674861
rect 563771 674593 563813 674829
rect 564049 674593 564091 674829
rect 563771 674509 564091 674593
rect 563771 674273 563813 674509
rect 564049 674273 564091 674509
rect 563771 674241 564091 674273
rect 573494 674829 574114 701273
rect 573494 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 574114 674829
rect 573494 674509 574114 674593
rect 573494 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 574114 674509
rect 22874 671454 23194 671486
rect 22874 671218 22916 671454
rect 23152 671218 23194 671454
rect 22874 671134 23194 671218
rect 22874 670898 22916 671134
rect 23152 670898 23194 671134
rect 22874 670866 23194 670898
rect 28805 671454 29125 671486
rect 28805 671218 28847 671454
rect 29083 671218 29125 671454
rect 28805 671134 29125 671218
rect 28805 670898 28847 671134
rect 29083 670898 29125 671134
rect 28805 670866 29125 670898
rect 50874 671454 51194 671486
rect 50874 671218 50916 671454
rect 51152 671218 51194 671454
rect 50874 671134 51194 671218
rect 50874 670898 50916 671134
rect 51152 670898 51194 671134
rect 50874 670866 51194 670898
rect 56805 671454 57125 671486
rect 56805 671218 56847 671454
rect 57083 671218 57125 671454
rect 56805 671134 57125 671218
rect 56805 670898 56847 671134
rect 57083 670898 57125 671134
rect 56805 670866 57125 670898
rect 78874 671454 79194 671486
rect 78874 671218 78916 671454
rect 79152 671218 79194 671454
rect 78874 671134 79194 671218
rect 78874 670898 78916 671134
rect 79152 670898 79194 671134
rect 78874 670866 79194 670898
rect 84805 671454 85125 671486
rect 84805 671218 84847 671454
rect 85083 671218 85125 671454
rect 84805 671134 85125 671218
rect 84805 670898 84847 671134
rect 85083 670898 85125 671134
rect 84805 670866 85125 670898
rect 106874 671454 107194 671486
rect 106874 671218 106916 671454
rect 107152 671218 107194 671454
rect 106874 671134 107194 671218
rect 106874 670898 106916 671134
rect 107152 670898 107194 671134
rect 106874 670866 107194 670898
rect 112805 671454 113125 671486
rect 112805 671218 112847 671454
rect 113083 671218 113125 671454
rect 112805 671134 113125 671218
rect 112805 670898 112847 671134
rect 113083 670898 113125 671134
rect 112805 670866 113125 670898
rect 134874 671454 135194 671486
rect 134874 671218 134916 671454
rect 135152 671218 135194 671454
rect 134874 671134 135194 671218
rect 134874 670898 134916 671134
rect 135152 670898 135194 671134
rect 134874 670866 135194 670898
rect 140805 671454 141125 671486
rect 140805 671218 140847 671454
rect 141083 671218 141125 671454
rect 140805 671134 141125 671218
rect 140805 670898 140847 671134
rect 141083 670898 141125 671134
rect 140805 670866 141125 670898
rect 162874 671454 163194 671486
rect 162874 671218 162916 671454
rect 163152 671218 163194 671454
rect 162874 671134 163194 671218
rect 162874 670898 162916 671134
rect 163152 670898 163194 671134
rect 162874 670866 163194 670898
rect 168805 671454 169125 671486
rect 168805 671218 168847 671454
rect 169083 671218 169125 671454
rect 168805 671134 169125 671218
rect 168805 670898 168847 671134
rect 169083 670898 169125 671134
rect 168805 670866 169125 670898
rect 190874 671454 191194 671486
rect 190874 671218 190916 671454
rect 191152 671218 191194 671454
rect 190874 671134 191194 671218
rect 190874 670898 190916 671134
rect 191152 670898 191194 671134
rect 190874 670866 191194 670898
rect 196805 671454 197125 671486
rect 196805 671218 196847 671454
rect 197083 671218 197125 671454
rect 196805 671134 197125 671218
rect 196805 670898 196847 671134
rect 197083 670898 197125 671134
rect 196805 670866 197125 670898
rect 218874 671454 219194 671486
rect 218874 671218 218916 671454
rect 219152 671218 219194 671454
rect 218874 671134 219194 671218
rect 218874 670898 218916 671134
rect 219152 670898 219194 671134
rect 218874 670866 219194 670898
rect 224805 671454 225125 671486
rect 224805 671218 224847 671454
rect 225083 671218 225125 671454
rect 224805 671134 225125 671218
rect 224805 670898 224847 671134
rect 225083 670898 225125 671134
rect 224805 670866 225125 670898
rect 246874 671454 247194 671486
rect 246874 671218 246916 671454
rect 247152 671218 247194 671454
rect 246874 671134 247194 671218
rect 246874 670898 246916 671134
rect 247152 670898 247194 671134
rect 246874 670866 247194 670898
rect 252805 671454 253125 671486
rect 252805 671218 252847 671454
rect 253083 671218 253125 671454
rect 252805 671134 253125 671218
rect 252805 670898 252847 671134
rect 253083 670898 253125 671134
rect 252805 670866 253125 670898
rect 274874 671454 275194 671486
rect 274874 671218 274916 671454
rect 275152 671218 275194 671454
rect 274874 671134 275194 671218
rect 274874 670898 274916 671134
rect 275152 670898 275194 671134
rect 274874 670866 275194 670898
rect 280805 671454 281125 671486
rect 280805 671218 280847 671454
rect 281083 671218 281125 671454
rect 280805 671134 281125 671218
rect 280805 670898 280847 671134
rect 281083 670898 281125 671134
rect 280805 670866 281125 670898
rect 302874 671454 303194 671486
rect 302874 671218 302916 671454
rect 303152 671218 303194 671454
rect 302874 671134 303194 671218
rect 302874 670898 302916 671134
rect 303152 670898 303194 671134
rect 302874 670866 303194 670898
rect 308805 671454 309125 671486
rect 308805 671218 308847 671454
rect 309083 671218 309125 671454
rect 308805 671134 309125 671218
rect 308805 670898 308847 671134
rect 309083 670898 309125 671134
rect 308805 670866 309125 670898
rect 330874 671454 331194 671486
rect 330874 671218 330916 671454
rect 331152 671218 331194 671454
rect 330874 671134 331194 671218
rect 330874 670898 330916 671134
rect 331152 670898 331194 671134
rect 330874 670866 331194 670898
rect 336805 671454 337125 671486
rect 336805 671218 336847 671454
rect 337083 671218 337125 671454
rect 336805 671134 337125 671218
rect 336805 670898 336847 671134
rect 337083 670898 337125 671134
rect 336805 670866 337125 670898
rect 358874 671454 359194 671486
rect 358874 671218 358916 671454
rect 359152 671218 359194 671454
rect 358874 671134 359194 671218
rect 358874 670898 358916 671134
rect 359152 670898 359194 671134
rect 358874 670866 359194 670898
rect 364805 671454 365125 671486
rect 364805 671218 364847 671454
rect 365083 671218 365125 671454
rect 364805 671134 365125 671218
rect 364805 670898 364847 671134
rect 365083 670898 365125 671134
rect 364805 670866 365125 670898
rect 386874 671454 387194 671486
rect 386874 671218 386916 671454
rect 387152 671218 387194 671454
rect 386874 671134 387194 671218
rect 386874 670898 386916 671134
rect 387152 670898 387194 671134
rect 386874 670866 387194 670898
rect 392805 671454 393125 671486
rect 392805 671218 392847 671454
rect 393083 671218 393125 671454
rect 392805 671134 393125 671218
rect 392805 670898 392847 671134
rect 393083 670898 393125 671134
rect 392805 670866 393125 670898
rect 414874 671454 415194 671486
rect 414874 671218 414916 671454
rect 415152 671218 415194 671454
rect 414874 671134 415194 671218
rect 414874 670898 414916 671134
rect 415152 670898 415194 671134
rect 414874 670866 415194 670898
rect 420805 671454 421125 671486
rect 420805 671218 420847 671454
rect 421083 671218 421125 671454
rect 420805 671134 421125 671218
rect 420805 670898 420847 671134
rect 421083 670898 421125 671134
rect 420805 670866 421125 670898
rect 442874 671454 443194 671486
rect 442874 671218 442916 671454
rect 443152 671218 443194 671454
rect 442874 671134 443194 671218
rect 442874 670898 442916 671134
rect 443152 670898 443194 671134
rect 442874 670866 443194 670898
rect 448805 671454 449125 671486
rect 448805 671218 448847 671454
rect 449083 671218 449125 671454
rect 448805 671134 449125 671218
rect 448805 670898 448847 671134
rect 449083 670898 449125 671134
rect 448805 670866 449125 670898
rect 470874 671454 471194 671486
rect 470874 671218 470916 671454
rect 471152 671218 471194 671454
rect 470874 671134 471194 671218
rect 470874 670898 470916 671134
rect 471152 670898 471194 671134
rect 470874 670866 471194 670898
rect 476805 671454 477125 671486
rect 476805 671218 476847 671454
rect 477083 671218 477125 671454
rect 476805 671134 477125 671218
rect 476805 670898 476847 671134
rect 477083 670898 477125 671134
rect 476805 670866 477125 670898
rect 498874 671454 499194 671486
rect 498874 671218 498916 671454
rect 499152 671218 499194 671454
rect 498874 671134 499194 671218
rect 498874 670898 498916 671134
rect 499152 670898 499194 671134
rect 498874 670866 499194 670898
rect 504805 671454 505125 671486
rect 504805 671218 504847 671454
rect 505083 671218 505125 671454
rect 504805 671134 505125 671218
rect 504805 670898 504847 671134
rect 505083 670898 505125 671134
rect 504805 670866 505125 670898
rect 526874 671454 527194 671486
rect 526874 671218 526916 671454
rect 527152 671218 527194 671454
rect 526874 671134 527194 671218
rect 526874 670898 526916 671134
rect 527152 670898 527194 671134
rect 526874 670866 527194 670898
rect 532805 671454 533125 671486
rect 532805 671218 532847 671454
rect 533083 671218 533125 671454
rect 532805 671134 533125 671218
rect 532805 670898 532847 671134
rect 533083 670898 533125 671134
rect 532805 670866 533125 670898
rect 554874 671454 555194 671486
rect 554874 671218 554916 671454
rect 555152 671218 555194 671454
rect 554874 671134 555194 671218
rect 554874 670898 554916 671134
rect 555152 670898 555194 671134
rect 554874 670866 555194 670898
rect 560805 671454 561125 671486
rect 560805 671218 560847 671454
rect 561083 671218 561125 671454
rect 560805 671134 561125 671218
rect 560805 670898 560847 671134
rect 561083 670898 561125 671134
rect 560805 670866 561125 670898
rect -2006 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 -1386 647829
rect -2006 647509 -1386 647593
rect -2006 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 -1386 647509
rect -2006 620829 -1386 647273
rect 19910 647829 20230 647861
rect 19910 647593 19952 647829
rect 20188 647593 20230 647829
rect 19910 647509 20230 647593
rect 19910 647273 19952 647509
rect 20188 647273 20230 647509
rect 19910 647241 20230 647273
rect 25840 647829 26160 647861
rect 25840 647593 25882 647829
rect 26118 647593 26160 647829
rect 25840 647509 26160 647593
rect 25840 647273 25882 647509
rect 26118 647273 26160 647509
rect 25840 647241 26160 647273
rect 31771 647829 32091 647861
rect 31771 647593 31813 647829
rect 32049 647593 32091 647829
rect 31771 647509 32091 647593
rect 31771 647273 31813 647509
rect 32049 647273 32091 647509
rect 31771 647241 32091 647273
rect 47910 647829 48230 647861
rect 47910 647593 47952 647829
rect 48188 647593 48230 647829
rect 47910 647509 48230 647593
rect 47910 647273 47952 647509
rect 48188 647273 48230 647509
rect 47910 647241 48230 647273
rect 53840 647829 54160 647861
rect 53840 647593 53882 647829
rect 54118 647593 54160 647829
rect 53840 647509 54160 647593
rect 53840 647273 53882 647509
rect 54118 647273 54160 647509
rect 53840 647241 54160 647273
rect 59771 647829 60091 647861
rect 59771 647593 59813 647829
rect 60049 647593 60091 647829
rect 59771 647509 60091 647593
rect 59771 647273 59813 647509
rect 60049 647273 60091 647509
rect 59771 647241 60091 647273
rect 75910 647829 76230 647861
rect 75910 647593 75952 647829
rect 76188 647593 76230 647829
rect 75910 647509 76230 647593
rect 75910 647273 75952 647509
rect 76188 647273 76230 647509
rect 75910 647241 76230 647273
rect 81840 647829 82160 647861
rect 81840 647593 81882 647829
rect 82118 647593 82160 647829
rect 81840 647509 82160 647593
rect 81840 647273 81882 647509
rect 82118 647273 82160 647509
rect 81840 647241 82160 647273
rect 87771 647829 88091 647861
rect 87771 647593 87813 647829
rect 88049 647593 88091 647829
rect 87771 647509 88091 647593
rect 87771 647273 87813 647509
rect 88049 647273 88091 647509
rect 87771 647241 88091 647273
rect 103910 647829 104230 647861
rect 103910 647593 103952 647829
rect 104188 647593 104230 647829
rect 103910 647509 104230 647593
rect 103910 647273 103952 647509
rect 104188 647273 104230 647509
rect 103910 647241 104230 647273
rect 109840 647829 110160 647861
rect 109840 647593 109882 647829
rect 110118 647593 110160 647829
rect 109840 647509 110160 647593
rect 109840 647273 109882 647509
rect 110118 647273 110160 647509
rect 109840 647241 110160 647273
rect 115771 647829 116091 647861
rect 115771 647593 115813 647829
rect 116049 647593 116091 647829
rect 115771 647509 116091 647593
rect 115771 647273 115813 647509
rect 116049 647273 116091 647509
rect 115771 647241 116091 647273
rect 131910 647829 132230 647861
rect 131910 647593 131952 647829
rect 132188 647593 132230 647829
rect 131910 647509 132230 647593
rect 131910 647273 131952 647509
rect 132188 647273 132230 647509
rect 131910 647241 132230 647273
rect 137840 647829 138160 647861
rect 137840 647593 137882 647829
rect 138118 647593 138160 647829
rect 137840 647509 138160 647593
rect 137840 647273 137882 647509
rect 138118 647273 138160 647509
rect 137840 647241 138160 647273
rect 143771 647829 144091 647861
rect 143771 647593 143813 647829
rect 144049 647593 144091 647829
rect 143771 647509 144091 647593
rect 143771 647273 143813 647509
rect 144049 647273 144091 647509
rect 143771 647241 144091 647273
rect 159910 647829 160230 647861
rect 159910 647593 159952 647829
rect 160188 647593 160230 647829
rect 159910 647509 160230 647593
rect 159910 647273 159952 647509
rect 160188 647273 160230 647509
rect 159910 647241 160230 647273
rect 165840 647829 166160 647861
rect 165840 647593 165882 647829
rect 166118 647593 166160 647829
rect 165840 647509 166160 647593
rect 165840 647273 165882 647509
rect 166118 647273 166160 647509
rect 165840 647241 166160 647273
rect 171771 647829 172091 647861
rect 171771 647593 171813 647829
rect 172049 647593 172091 647829
rect 171771 647509 172091 647593
rect 171771 647273 171813 647509
rect 172049 647273 172091 647509
rect 171771 647241 172091 647273
rect 187910 647829 188230 647861
rect 187910 647593 187952 647829
rect 188188 647593 188230 647829
rect 187910 647509 188230 647593
rect 187910 647273 187952 647509
rect 188188 647273 188230 647509
rect 187910 647241 188230 647273
rect 193840 647829 194160 647861
rect 193840 647593 193882 647829
rect 194118 647593 194160 647829
rect 193840 647509 194160 647593
rect 193840 647273 193882 647509
rect 194118 647273 194160 647509
rect 193840 647241 194160 647273
rect 199771 647829 200091 647861
rect 199771 647593 199813 647829
rect 200049 647593 200091 647829
rect 199771 647509 200091 647593
rect 199771 647273 199813 647509
rect 200049 647273 200091 647509
rect 199771 647241 200091 647273
rect 215910 647829 216230 647861
rect 215910 647593 215952 647829
rect 216188 647593 216230 647829
rect 215910 647509 216230 647593
rect 215910 647273 215952 647509
rect 216188 647273 216230 647509
rect 215910 647241 216230 647273
rect 221840 647829 222160 647861
rect 221840 647593 221882 647829
rect 222118 647593 222160 647829
rect 221840 647509 222160 647593
rect 221840 647273 221882 647509
rect 222118 647273 222160 647509
rect 221840 647241 222160 647273
rect 227771 647829 228091 647861
rect 227771 647593 227813 647829
rect 228049 647593 228091 647829
rect 227771 647509 228091 647593
rect 227771 647273 227813 647509
rect 228049 647273 228091 647509
rect 227771 647241 228091 647273
rect 243910 647829 244230 647861
rect 243910 647593 243952 647829
rect 244188 647593 244230 647829
rect 243910 647509 244230 647593
rect 243910 647273 243952 647509
rect 244188 647273 244230 647509
rect 243910 647241 244230 647273
rect 249840 647829 250160 647861
rect 249840 647593 249882 647829
rect 250118 647593 250160 647829
rect 249840 647509 250160 647593
rect 249840 647273 249882 647509
rect 250118 647273 250160 647509
rect 249840 647241 250160 647273
rect 255771 647829 256091 647861
rect 255771 647593 255813 647829
rect 256049 647593 256091 647829
rect 255771 647509 256091 647593
rect 255771 647273 255813 647509
rect 256049 647273 256091 647509
rect 255771 647241 256091 647273
rect 271910 647829 272230 647861
rect 271910 647593 271952 647829
rect 272188 647593 272230 647829
rect 271910 647509 272230 647593
rect 271910 647273 271952 647509
rect 272188 647273 272230 647509
rect 271910 647241 272230 647273
rect 277840 647829 278160 647861
rect 277840 647593 277882 647829
rect 278118 647593 278160 647829
rect 277840 647509 278160 647593
rect 277840 647273 277882 647509
rect 278118 647273 278160 647509
rect 277840 647241 278160 647273
rect 283771 647829 284091 647861
rect 283771 647593 283813 647829
rect 284049 647593 284091 647829
rect 283771 647509 284091 647593
rect 283771 647273 283813 647509
rect 284049 647273 284091 647509
rect 283771 647241 284091 647273
rect 299910 647829 300230 647861
rect 299910 647593 299952 647829
rect 300188 647593 300230 647829
rect 299910 647509 300230 647593
rect 299910 647273 299952 647509
rect 300188 647273 300230 647509
rect 299910 647241 300230 647273
rect 305840 647829 306160 647861
rect 305840 647593 305882 647829
rect 306118 647593 306160 647829
rect 305840 647509 306160 647593
rect 305840 647273 305882 647509
rect 306118 647273 306160 647509
rect 305840 647241 306160 647273
rect 311771 647829 312091 647861
rect 311771 647593 311813 647829
rect 312049 647593 312091 647829
rect 311771 647509 312091 647593
rect 311771 647273 311813 647509
rect 312049 647273 312091 647509
rect 311771 647241 312091 647273
rect 327910 647829 328230 647861
rect 327910 647593 327952 647829
rect 328188 647593 328230 647829
rect 327910 647509 328230 647593
rect 327910 647273 327952 647509
rect 328188 647273 328230 647509
rect 327910 647241 328230 647273
rect 333840 647829 334160 647861
rect 333840 647593 333882 647829
rect 334118 647593 334160 647829
rect 333840 647509 334160 647593
rect 333840 647273 333882 647509
rect 334118 647273 334160 647509
rect 333840 647241 334160 647273
rect 339771 647829 340091 647861
rect 339771 647593 339813 647829
rect 340049 647593 340091 647829
rect 339771 647509 340091 647593
rect 339771 647273 339813 647509
rect 340049 647273 340091 647509
rect 339771 647241 340091 647273
rect 355910 647829 356230 647861
rect 355910 647593 355952 647829
rect 356188 647593 356230 647829
rect 355910 647509 356230 647593
rect 355910 647273 355952 647509
rect 356188 647273 356230 647509
rect 355910 647241 356230 647273
rect 361840 647829 362160 647861
rect 361840 647593 361882 647829
rect 362118 647593 362160 647829
rect 361840 647509 362160 647593
rect 361840 647273 361882 647509
rect 362118 647273 362160 647509
rect 361840 647241 362160 647273
rect 367771 647829 368091 647861
rect 367771 647593 367813 647829
rect 368049 647593 368091 647829
rect 367771 647509 368091 647593
rect 367771 647273 367813 647509
rect 368049 647273 368091 647509
rect 367771 647241 368091 647273
rect 383910 647829 384230 647861
rect 383910 647593 383952 647829
rect 384188 647593 384230 647829
rect 383910 647509 384230 647593
rect 383910 647273 383952 647509
rect 384188 647273 384230 647509
rect 383910 647241 384230 647273
rect 389840 647829 390160 647861
rect 389840 647593 389882 647829
rect 390118 647593 390160 647829
rect 389840 647509 390160 647593
rect 389840 647273 389882 647509
rect 390118 647273 390160 647509
rect 389840 647241 390160 647273
rect 395771 647829 396091 647861
rect 395771 647593 395813 647829
rect 396049 647593 396091 647829
rect 395771 647509 396091 647593
rect 395771 647273 395813 647509
rect 396049 647273 396091 647509
rect 395771 647241 396091 647273
rect 411910 647829 412230 647861
rect 411910 647593 411952 647829
rect 412188 647593 412230 647829
rect 411910 647509 412230 647593
rect 411910 647273 411952 647509
rect 412188 647273 412230 647509
rect 411910 647241 412230 647273
rect 417840 647829 418160 647861
rect 417840 647593 417882 647829
rect 418118 647593 418160 647829
rect 417840 647509 418160 647593
rect 417840 647273 417882 647509
rect 418118 647273 418160 647509
rect 417840 647241 418160 647273
rect 423771 647829 424091 647861
rect 423771 647593 423813 647829
rect 424049 647593 424091 647829
rect 423771 647509 424091 647593
rect 423771 647273 423813 647509
rect 424049 647273 424091 647509
rect 423771 647241 424091 647273
rect 439910 647829 440230 647861
rect 439910 647593 439952 647829
rect 440188 647593 440230 647829
rect 439910 647509 440230 647593
rect 439910 647273 439952 647509
rect 440188 647273 440230 647509
rect 439910 647241 440230 647273
rect 445840 647829 446160 647861
rect 445840 647593 445882 647829
rect 446118 647593 446160 647829
rect 445840 647509 446160 647593
rect 445840 647273 445882 647509
rect 446118 647273 446160 647509
rect 445840 647241 446160 647273
rect 451771 647829 452091 647861
rect 451771 647593 451813 647829
rect 452049 647593 452091 647829
rect 451771 647509 452091 647593
rect 451771 647273 451813 647509
rect 452049 647273 452091 647509
rect 451771 647241 452091 647273
rect 467910 647829 468230 647861
rect 467910 647593 467952 647829
rect 468188 647593 468230 647829
rect 467910 647509 468230 647593
rect 467910 647273 467952 647509
rect 468188 647273 468230 647509
rect 467910 647241 468230 647273
rect 473840 647829 474160 647861
rect 473840 647593 473882 647829
rect 474118 647593 474160 647829
rect 473840 647509 474160 647593
rect 473840 647273 473882 647509
rect 474118 647273 474160 647509
rect 473840 647241 474160 647273
rect 479771 647829 480091 647861
rect 479771 647593 479813 647829
rect 480049 647593 480091 647829
rect 479771 647509 480091 647593
rect 479771 647273 479813 647509
rect 480049 647273 480091 647509
rect 479771 647241 480091 647273
rect 495910 647829 496230 647861
rect 495910 647593 495952 647829
rect 496188 647593 496230 647829
rect 495910 647509 496230 647593
rect 495910 647273 495952 647509
rect 496188 647273 496230 647509
rect 495910 647241 496230 647273
rect 501840 647829 502160 647861
rect 501840 647593 501882 647829
rect 502118 647593 502160 647829
rect 501840 647509 502160 647593
rect 501840 647273 501882 647509
rect 502118 647273 502160 647509
rect 501840 647241 502160 647273
rect 507771 647829 508091 647861
rect 507771 647593 507813 647829
rect 508049 647593 508091 647829
rect 507771 647509 508091 647593
rect 507771 647273 507813 647509
rect 508049 647273 508091 647509
rect 507771 647241 508091 647273
rect 523910 647829 524230 647861
rect 523910 647593 523952 647829
rect 524188 647593 524230 647829
rect 523910 647509 524230 647593
rect 523910 647273 523952 647509
rect 524188 647273 524230 647509
rect 523910 647241 524230 647273
rect 529840 647829 530160 647861
rect 529840 647593 529882 647829
rect 530118 647593 530160 647829
rect 529840 647509 530160 647593
rect 529840 647273 529882 647509
rect 530118 647273 530160 647509
rect 529840 647241 530160 647273
rect 535771 647829 536091 647861
rect 535771 647593 535813 647829
rect 536049 647593 536091 647829
rect 535771 647509 536091 647593
rect 535771 647273 535813 647509
rect 536049 647273 536091 647509
rect 535771 647241 536091 647273
rect 551910 647829 552230 647861
rect 551910 647593 551952 647829
rect 552188 647593 552230 647829
rect 551910 647509 552230 647593
rect 551910 647273 551952 647509
rect 552188 647273 552230 647509
rect 551910 647241 552230 647273
rect 557840 647829 558160 647861
rect 557840 647593 557882 647829
rect 558118 647593 558160 647829
rect 557840 647509 558160 647593
rect 557840 647273 557882 647509
rect 558118 647273 558160 647509
rect 557840 647241 558160 647273
rect 563771 647829 564091 647861
rect 563771 647593 563813 647829
rect 564049 647593 564091 647829
rect 563771 647509 564091 647593
rect 563771 647273 563813 647509
rect 564049 647273 564091 647509
rect 563771 647241 564091 647273
rect 573494 647829 574114 674273
rect 573494 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 574114 647829
rect 573494 647509 574114 647593
rect 573494 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 574114 647509
rect 22874 644454 23194 644486
rect 22874 644218 22916 644454
rect 23152 644218 23194 644454
rect 22874 644134 23194 644218
rect 22874 643898 22916 644134
rect 23152 643898 23194 644134
rect 22874 643866 23194 643898
rect 28805 644454 29125 644486
rect 28805 644218 28847 644454
rect 29083 644218 29125 644454
rect 28805 644134 29125 644218
rect 28805 643898 28847 644134
rect 29083 643898 29125 644134
rect 28805 643866 29125 643898
rect 50874 644454 51194 644486
rect 50874 644218 50916 644454
rect 51152 644218 51194 644454
rect 50874 644134 51194 644218
rect 50874 643898 50916 644134
rect 51152 643898 51194 644134
rect 50874 643866 51194 643898
rect 56805 644454 57125 644486
rect 56805 644218 56847 644454
rect 57083 644218 57125 644454
rect 56805 644134 57125 644218
rect 56805 643898 56847 644134
rect 57083 643898 57125 644134
rect 56805 643866 57125 643898
rect 78874 644454 79194 644486
rect 78874 644218 78916 644454
rect 79152 644218 79194 644454
rect 78874 644134 79194 644218
rect 78874 643898 78916 644134
rect 79152 643898 79194 644134
rect 78874 643866 79194 643898
rect 84805 644454 85125 644486
rect 84805 644218 84847 644454
rect 85083 644218 85125 644454
rect 84805 644134 85125 644218
rect 84805 643898 84847 644134
rect 85083 643898 85125 644134
rect 84805 643866 85125 643898
rect 106874 644454 107194 644486
rect 106874 644218 106916 644454
rect 107152 644218 107194 644454
rect 106874 644134 107194 644218
rect 106874 643898 106916 644134
rect 107152 643898 107194 644134
rect 106874 643866 107194 643898
rect 112805 644454 113125 644486
rect 112805 644218 112847 644454
rect 113083 644218 113125 644454
rect 112805 644134 113125 644218
rect 112805 643898 112847 644134
rect 113083 643898 113125 644134
rect 112805 643866 113125 643898
rect 134874 644454 135194 644486
rect 134874 644218 134916 644454
rect 135152 644218 135194 644454
rect 134874 644134 135194 644218
rect 134874 643898 134916 644134
rect 135152 643898 135194 644134
rect 134874 643866 135194 643898
rect 140805 644454 141125 644486
rect 140805 644218 140847 644454
rect 141083 644218 141125 644454
rect 140805 644134 141125 644218
rect 140805 643898 140847 644134
rect 141083 643898 141125 644134
rect 140805 643866 141125 643898
rect 162874 644454 163194 644486
rect 162874 644218 162916 644454
rect 163152 644218 163194 644454
rect 162874 644134 163194 644218
rect 162874 643898 162916 644134
rect 163152 643898 163194 644134
rect 162874 643866 163194 643898
rect 168805 644454 169125 644486
rect 168805 644218 168847 644454
rect 169083 644218 169125 644454
rect 168805 644134 169125 644218
rect 168805 643898 168847 644134
rect 169083 643898 169125 644134
rect 168805 643866 169125 643898
rect 190874 644454 191194 644486
rect 190874 644218 190916 644454
rect 191152 644218 191194 644454
rect 190874 644134 191194 644218
rect 190874 643898 190916 644134
rect 191152 643898 191194 644134
rect 190874 643866 191194 643898
rect 196805 644454 197125 644486
rect 196805 644218 196847 644454
rect 197083 644218 197125 644454
rect 196805 644134 197125 644218
rect 196805 643898 196847 644134
rect 197083 643898 197125 644134
rect 196805 643866 197125 643898
rect 218874 644454 219194 644486
rect 218874 644218 218916 644454
rect 219152 644218 219194 644454
rect 218874 644134 219194 644218
rect 218874 643898 218916 644134
rect 219152 643898 219194 644134
rect 218874 643866 219194 643898
rect 224805 644454 225125 644486
rect 224805 644218 224847 644454
rect 225083 644218 225125 644454
rect 224805 644134 225125 644218
rect 224805 643898 224847 644134
rect 225083 643898 225125 644134
rect 224805 643866 225125 643898
rect 246874 644454 247194 644486
rect 246874 644218 246916 644454
rect 247152 644218 247194 644454
rect 246874 644134 247194 644218
rect 246874 643898 246916 644134
rect 247152 643898 247194 644134
rect 246874 643866 247194 643898
rect 252805 644454 253125 644486
rect 252805 644218 252847 644454
rect 253083 644218 253125 644454
rect 252805 644134 253125 644218
rect 252805 643898 252847 644134
rect 253083 643898 253125 644134
rect 252805 643866 253125 643898
rect 274874 644454 275194 644486
rect 274874 644218 274916 644454
rect 275152 644218 275194 644454
rect 274874 644134 275194 644218
rect 274874 643898 274916 644134
rect 275152 643898 275194 644134
rect 274874 643866 275194 643898
rect 280805 644454 281125 644486
rect 280805 644218 280847 644454
rect 281083 644218 281125 644454
rect 280805 644134 281125 644218
rect 280805 643898 280847 644134
rect 281083 643898 281125 644134
rect 280805 643866 281125 643898
rect 302874 644454 303194 644486
rect 302874 644218 302916 644454
rect 303152 644218 303194 644454
rect 302874 644134 303194 644218
rect 302874 643898 302916 644134
rect 303152 643898 303194 644134
rect 302874 643866 303194 643898
rect 308805 644454 309125 644486
rect 308805 644218 308847 644454
rect 309083 644218 309125 644454
rect 308805 644134 309125 644218
rect 308805 643898 308847 644134
rect 309083 643898 309125 644134
rect 308805 643866 309125 643898
rect 330874 644454 331194 644486
rect 330874 644218 330916 644454
rect 331152 644218 331194 644454
rect 330874 644134 331194 644218
rect 330874 643898 330916 644134
rect 331152 643898 331194 644134
rect 330874 643866 331194 643898
rect 336805 644454 337125 644486
rect 336805 644218 336847 644454
rect 337083 644218 337125 644454
rect 336805 644134 337125 644218
rect 336805 643898 336847 644134
rect 337083 643898 337125 644134
rect 336805 643866 337125 643898
rect 358874 644454 359194 644486
rect 358874 644218 358916 644454
rect 359152 644218 359194 644454
rect 358874 644134 359194 644218
rect 358874 643898 358916 644134
rect 359152 643898 359194 644134
rect 358874 643866 359194 643898
rect 364805 644454 365125 644486
rect 364805 644218 364847 644454
rect 365083 644218 365125 644454
rect 364805 644134 365125 644218
rect 364805 643898 364847 644134
rect 365083 643898 365125 644134
rect 364805 643866 365125 643898
rect 386874 644454 387194 644486
rect 386874 644218 386916 644454
rect 387152 644218 387194 644454
rect 386874 644134 387194 644218
rect 386874 643898 386916 644134
rect 387152 643898 387194 644134
rect 386874 643866 387194 643898
rect 392805 644454 393125 644486
rect 392805 644218 392847 644454
rect 393083 644218 393125 644454
rect 392805 644134 393125 644218
rect 392805 643898 392847 644134
rect 393083 643898 393125 644134
rect 392805 643866 393125 643898
rect 414874 644454 415194 644486
rect 414874 644218 414916 644454
rect 415152 644218 415194 644454
rect 414874 644134 415194 644218
rect 414874 643898 414916 644134
rect 415152 643898 415194 644134
rect 414874 643866 415194 643898
rect 420805 644454 421125 644486
rect 420805 644218 420847 644454
rect 421083 644218 421125 644454
rect 420805 644134 421125 644218
rect 420805 643898 420847 644134
rect 421083 643898 421125 644134
rect 420805 643866 421125 643898
rect 442874 644454 443194 644486
rect 442874 644218 442916 644454
rect 443152 644218 443194 644454
rect 442874 644134 443194 644218
rect 442874 643898 442916 644134
rect 443152 643898 443194 644134
rect 442874 643866 443194 643898
rect 448805 644454 449125 644486
rect 448805 644218 448847 644454
rect 449083 644218 449125 644454
rect 448805 644134 449125 644218
rect 448805 643898 448847 644134
rect 449083 643898 449125 644134
rect 448805 643866 449125 643898
rect 470874 644454 471194 644486
rect 470874 644218 470916 644454
rect 471152 644218 471194 644454
rect 470874 644134 471194 644218
rect 470874 643898 470916 644134
rect 471152 643898 471194 644134
rect 470874 643866 471194 643898
rect 476805 644454 477125 644486
rect 476805 644218 476847 644454
rect 477083 644218 477125 644454
rect 476805 644134 477125 644218
rect 476805 643898 476847 644134
rect 477083 643898 477125 644134
rect 476805 643866 477125 643898
rect 498874 644454 499194 644486
rect 498874 644218 498916 644454
rect 499152 644218 499194 644454
rect 498874 644134 499194 644218
rect 498874 643898 498916 644134
rect 499152 643898 499194 644134
rect 498874 643866 499194 643898
rect 504805 644454 505125 644486
rect 504805 644218 504847 644454
rect 505083 644218 505125 644454
rect 504805 644134 505125 644218
rect 504805 643898 504847 644134
rect 505083 643898 505125 644134
rect 504805 643866 505125 643898
rect 526874 644454 527194 644486
rect 526874 644218 526916 644454
rect 527152 644218 527194 644454
rect 526874 644134 527194 644218
rect 526874 643898 526916 644134
rect 527152 643898 527194 644134
rect 526874 643866 527194 643898
rect 532805 644454 533125 644486
rect 532805 644218 532847 644454
rect 533083 644218 533125 644454
rect 532805 644134 533125 644218
rect 532805 643898 532847 644134
rect 533083 643898 533125 644134
rect 532805 643866 533125 643898
rect 554874 644454 555194 644486
rect 554874 644218 554916 644454
rect 555152 644218 555194 644454
rect 554874 644134 555194 644218
rect 554874 643898 554916 644134
rect 555152 643898 555194 644134
rect 554874 643866 555194 643898
rect 560805 644454 561125 644486
rect 560805 644218 560847 644454
rect 561083 644218 561125 644454
rect 560805 644134 561125 644218
rect 560805 643898 560847 644134
rect 561083 643898 561125 644134
rect 560805 643866 561125 643898
rect -2006 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 -1386 620829
rect -2006 620509 -1386 620593
rect -2006 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 -1386 620509
rect -2006 593829 -1386 620273
rect 19910 620829 20230 620861
rect 19910 620593 19952 620829
rect 20188 620593 20230 620829
rect 19910 620509 20230 620593
rect 19910 620273 19952 620509
rect 20188 620273 20230 620509
rect 19910 620241 20230 620273
rect 25840 620829 26160 620861
rect 25840 620593 25882 620829
rect 26118 620593 26160 620829
rect 25840 620509 26160 620593
rect 25840 620273 25882 620509
rect 26118 620273 26160 620509
rect 25840 620241 26160 620273
rect 31771 620829 32091 620861
rect 31771 620593 31813 620829
rect 32049 620593 32091 620829
rect 31771 620509 32091 620593
rect 31771 620273 31813 620509
rect 32049 620273 32091 620509
rect 31771 620241 32091 620273
rect 47910 620829 48230 620861
rect 47910 620593 47952 620829
rect 48188 620593 48230 620829
rect 47910 620509 48230 620593
rect 47910 620273 47952 620509
rect 48188 620273 48230 620509
rect 47910 620241 48230 620273
rect 53840 620829 54160 620861
rect 53840 620593 53882 620829
rect 54118 620593 54160 620829
rect 53840 620509 54160 620593
rect 53840 620273 53882 620509
rect 54118 620273 54160 620509
rect 53840 620241 54160 620273
rect 59771 620829 60091 620861
rect 59771 620593 59813 620829
rect 60049 620593 60091 620829
rect 59771 620509 60091 620593
rect 59771 620273 59813 620509
rect 60049 620273 60091 620509
rect 59771 620241 60091 620273
rect 75910 620829 76230 620861
rect 75910 620593 75952 620829
rect 76188 620593 76230 620829
rect 75910 620509 76230 620593
rect 75910 620273 75952 620509
rect 76188 620273 76230 620509
rect 75910 620241 76230 620273
rect 81840 620829 82160 620861
rect 81840 620593 81882 620829
rect 82118 620593 82160 620829
rect 81840 620509 82160 620593
rect 81840 620273 81882 620509
rect 82118 620273 82160 620509
rect 81840 620241 82160 620273
rect 87771 620829 88091 620861
rect 87771 620593 87813 620829
rect 88049 620593 88091 620829
rect 87771 620509 88091 620593
rect 87771 620273 87813 620509
rect 88049 620273 88091 620509
rect 87771 620241 88091 620273
rect 103910 620829 104230 620861
rect 103910 620593 103952 620829
rect 104188 620593 104230 620829
rect 103910 620509 104230 620593
rect 103910 620273 103952 620509
rect 104188 620273 104230 620509
rect 103910 620241 104230 620273
rect 109840 620829 110160 620861
rect 109840 620593 109882 620829
rect 110118 620593 110160 620829
rect 109840 620509 110160 620593
rect 109840 620273 109882 620509
rect 110118 620273 110160 620509
rect 109840 620241 110160 620273
rect 115771 620829 116091 620861
rect 115771 620593 115813 620829
rect 116049 620593 116091 620829
rect 115771 620509 116091 620593
rect 115771 620273 115813 620509
rect 116049 620273 116091 620509
rect 115771 620241 116091 620273
rect 131910 620829 132230 620861
rect 131910 620593 131952 620829
rect 132188 620593 132230 620829
rect 131910 620509 132230 620593
rect 131910 620273 131952 620509
rect 132188 620273 132230 620509
rect 131910 620241 132230 620273
rect 137840 620829 138160 620861
rect 137840 620593 137882 620829
rect 138118 620593 138160 620829
rect 137840 620509 138160 620593
rect 137840 620273 137882 620509
rect 138118 620273 138160 620509
rect 137840 620241 138160 620273
rect 143771 620829 144091 620861
rect 143771 620593 143813 620829
rect 144049 620593 144091 620829
rect 143771 620509 144091 620593
rect 143771 620273 143813 620509
rect 144049 620273 144091 620509
rect 143771 620241 144091 620273
rect 159910 620829 160230 620861
rect 159910 620593 159952 620829
rect 160188 620593 160230 620829
rect 159910 620509 160230 620593
rect 159910 620273 159952 620509
rect 160188 620273 160230 620509
rect 159910 620241 160230 620273
rect 165840 620829 166160 620861
rect 165840 620593 165882 620829
rect 166118 620593 166160 620829
rect 165840 620509 166160 620593
rect 165840 620273 165882 620509
rect 166118 620273 166160 620509
rect 165840 620241 166160 620273
rect 171771 620829 172091 620861
rect 171771 620593 171813 620829
rect 172049 620593 172091 620829
rect 171771 620509 172091 620593
rect 171771 620273 171813 620509
rect 172049 620273 172091 620509
rect 171771 620241 172091 620273
rect 187910 620829 188230 620861
rect 187910 620593 187952 620829
rect 188188 620593 188230 620829
rect 187910 620509 188230 620593
rect 187910 620273 187952 620509
rect 188188 620273 188230 620509
rect 187910 620241 188230 620273
rect 193840 620829 194160 620861
rect 193840 620593 193882 620829
rect 194118 620593 194160 620829
rect 193840 620509 194160 620593
rect 193840 620273 193882 620509
rect 194118 620273 194160 620509
rect 193840 620241 194160 620273
rect 199771 620829 200091 620861
rect 199771 620593 199813 620829
rect 200049 620593 200091 620829
rect 199771 620509 200091 620593
rect 199771 620273 199813 620509
rect 200049 620273 200091 620509
rect 199771 620241 200091 620273
rect 215910 620829 216230 620861
rect 215910 620593 215952 620829
rect 216188 620593 216230 620829
rect 215910 620509 216230 620593
rect 215910 620273 215952 620509
rect 216188 620273 216230 620509
rect 215910 620241 216230 620273
rect 221840 620829 222160 620861
rect 221840 620593 221882 620829
rect 222118 620593 222160 620829
rect 221840 620509 222160 620593
rect 221840 620273 221882 620509
rect 222118 620273 222160 620509
rect 221840 620241 222160 620273
rect 227771 620829 228091 620861
rect 227771 620593 227813 620829
rect 228049 620593 228091 620829
rect 227771 620509 228091 620593
rect 227771 620273 227813 620509
rect 228049 620273 228091 620509
rect 227771 620241 228091 620273
rect 243910 620829 244230 620861
rect 243910 620593 243952 620829
rect 244188 620593 244230 620829
rect 243910 620509 244230 620593
rect 243910 620273 243952 620509
rect 244188 620273 244230 620509
rect 243910 620241 244230 620273
rect 249840 620829 250160 620861
rect 249840 620593 249882 620829
rect 250118 620593 250160 620829
rect 249840 620509 250160 620593
rect 249840 620273 249882 620509
rect 250118 620273 250160 620509
rect 249840 620241 250160 620273
rect 255771 620829 256091 620861
rect 255771 620593 255813 620829
rect 256049 620593 256091 620829
rect 255771 620509 256091 620593
rect 255771 620273 255813 620509
rect 256049 620273 256091 620509
rect 255771 620241 256091 620273
rect 271910 620829 272230 620861
rect 271910 620593 271952 620829
rect 272188 620593 272230 620829
rect 271910 620509 272230 620593
rect 271910 620273 271952 620509
rect 272188 620273 272230 620509
rect 271910 620241 272230 620273
rect 277840 620829 278160 620861
rect 277840 620593 277882 620829
rect 278118 620593 278160 620829
rect 277840 620509 278160 620593
rect 277840 620273 277882 620509
rect 278118 620273 278160 620509
rect 277840 620241 278160 620273
rect 283771 620829 284091 620861
rect 283771 620593 283813 620829
rect 284049 620593 284091 620829
rect 283771 620509 284091 620593
rect 283771 620273 283813 620509
rect 284049 620273 284091 620509
rect 283771 620241 284091 620273
rect 299910 620829 300230 620861
rect 299910 620593 299952 620829
rect 300188 620593 300230 620829
rect 299910 620509 300230 620593
rect 299910 620273 299952 620509
rect 300188 620273 300230 620509
rect 299910 620241 300230 620273
rect 305840 620829 306160 620861
rect 305840 620593 305882 620829
rect 306118 620593 306160 620829
rect 305840 620509 306160 620593
rect 305840 620273 305882 620509
rect 306118 620273 306160 620509
rect 305840 620241 306160 620273
rect 311771 620829 312091 620861
rect 311771 620593 311813 620829
rect 312049 620593 312091 620829
rect 311771 620509 312091 620593
rect 311771 620273 311813 620509
rect 312049 620273 312091 620509
rect 311771 620241 312091 620273
rect 327910 620829 328230 620861
rect 327910 620593 327952 620829
rect 328188 620593 328230 620829
rect 327910 620509 328230 620593
rect 327910 620273 327952 620509
rect 328188 620273 328230 620509
rect 327910 620241 328230 620273
rect 333840 620829 334160 620861
rect 333840 620593 333882 620829
rect 334118 620593 334160 620829
rect 333840 620509 334160 620593
rect 333840 620273 333882 620509
rect 334118 620273 334160 620509
rect 333840 620241 334160 620273
rect 339771 620829 340091 620861
rect 339771 620593 339813 620829
rect 340049 620593 340091 620829
rect 339771 620509 340091 620593
rect 339771 620273 339813 620509
rect 340049 620273 340091 620509
rect 339771 620241 340091 620273
rect 355910 620829 356230 620861
rect 355910 620593 355952 620829
rect 356188 620593 356230 620829
rect 355910 620509 356230 620593
rect 355910 620273 355952 620509
rect 356188 620273 356230 620509
rect 355910 620241 356230 620273
rect 361840 620829 362160 620861
rect 361840 620593 361882 620829
rect 362118 620593 362160 620829
rect 361840 620509 362160 620593
rect 361840 620273 361882 620509
rect 362118 620273 362160 620509
rect 361840 620241 362160 620273
rect 367771 620829 368091 620861
rect 367771 620593 367813 620829
rect 368049 620593 368091 620829
rect 367771 620509 368091 620593
rect 367771 620273 367813 620509
rect 368049 620273 368091 620509
rect 367771 620241 368091 620273
rect 383910 620829 384230 620861
rect 383910 620593 383952 620829
rect 384188 620593 384230 620829
rect 383910 620509 384230 620593
rect 383910 620273 383952 620509
rect 384188 620273 384230 620509
rect 383910 620241 384230 620273
rect 389840 620829 390160 620861
rect 389840 620593 389882 620829
rect 390118 620593 390160 620829
rect 389840 620509 390160 620593
rect 389840 620273 389882 620509
rect 390118 620273 390160 620509
rect 389840 620241 390160 620273
rect 395771 620829 396091 620861
rect 395771 620593 395813 620829
rect 396049 620593 396091 620829
rect 395771 620509 396091 620593
rect 395771 620273 395813 620509
rect 396049 620273 396091 620509
rect 395771 620241 396091 620273
rect 411910 620829 412230 620861
rect 411910 620593 411952 620829
rect 412188 620593 412230 620829
rect 411910 620509 412230 620593
rect 411910 620273 411952 620509
rect 412188 620273 412230 620509
rect 411910 620241 412230 620273
rect 417840 620829 418160 620861
rect 417840 620593 417882 620829
rect 418118 620593 418160 620829
rect 417840 620509 418160 620593
rect 417840 620273 417882 620509
rect 418118 620273 418160 620509
rect 417840 620241 418160 620273
rect 423771 620829 424091 620861
rect 423771 620593 423813 620829
rect 424049 620593 424091 620829
rect 423771 620509 424091 620593
rect 423771 620273 423813 620509
rect 424049 620273 424091 620509
rect 423771 620241 424091 620273
rect 439910 620829 440230 620861
rect 439910 620593 439952 620829
rect 440188 620593 440230 620829
rect 439910 620509 440230 620593
rect 439910 620273 439952 620509
rect 440188 620273 440230 620509
rect 439910 620241 440230 620273
rect 445840 620829 446160 620861
rect 445840 620593 445882 620829
rect 446118 620593 446160 620829
rect 445840 620509 446160 620593
rect 445840 620273 445882 620509
rect 446118 620273 446160 620509
rect 445840 620241 446160 620273
rect 451771 620829 452091 620861
rect 451771 620593 451813 620829
rect 452049 620593 452091 620829
rect 451771 620509 452091 620593
rect 451771 620273 451813 620509
rect 452049 620273 452091 620509
rect 451771 620241 452091 620273
rect 467910 620829 468230 620861
rect 467910 620593 467952 620829
rect 468188 620593 468230 620829
rect 467910 620509 468230 620593
rect 467910 620273 467952 620509
rect 468188 620273 468230 620509
rect 467910 620241 468230 620273
rect 473840 620829 474160 620861
rect 473840 620593 473882 620829
rect 474118 620593 474160 620829
rect 473840 620509 474160 620593
rect 473840 620273 473882 620509
rect 474118 620273 474160 620509
rect 473840 620241 474160 620273
rect 479771 620829 480091 620861
rect 479771 620593 479813 620829
rect 480049 620593 480091 620829
rect 479771 620509 480091 620593
rect 479771 620273 479813 620509
rect 480049 620273 480091 620509
rect 479771 620241 480091 620273
rect 495910 620829 496230 620861
rect 495910 620593 495952 620829
rect 496188 620593 496230 620829
rect 495910 620509 496230 620593
rect 495910 620273 495952 620509
rect 496188 620273 496230 620509
rect 495910 620241 496230 620273
rect 501840 620829 502160 620861
rect 501840 620593 501882 620829
rect 502118 620593 502160 620829
rect 501840 620509 502160 620593
rect 501840 620273 501882 620509
rect 502118 620273 502160 620509
rect 501840 620241 502160 620273
rect 507771 620829 508091 620861
rect 507771 620593 507813 620829
rect 508049 620593 508091 620829
rect 507771 620509 508091 620593
rect 507771 620273 507813 620509
rect 508049 620273 508091 620509
rect 507771 620241 508091 620273
rect 523910 620829 524230 620861
rect 523910 620593 523952 620829
rect 524188 620593 524230 620829
rect 523910 620509 524230 620593
rect 523910 620273 523952 620509
rect 524188 620273 524230 620509
rect 523910 620241 524230 620273
rect 529840 620829 530160 620861
rect 529840 620593 529882 620829
rect 530118 620593 530160 620829
rect 529840 620509 530160 620593
rect 529840 620273 529882 620509
rect 530118 620273 530160 620509
rect 529840 620241 530160 620273
rect 535771 620829 536091 620861
rect 535771 620593 535813 620829
rect 536049 620593 536091 620829
rect 535771 620509 536091 620593
rect 535771 620273 535813 620509
rect 536049 620273 536091 620509
rect 535771 620241 536091 620273
rect 551910 620829 552230 620861
rect 551910 620593 551952 620829
rect 552188 620593 552230 620829
rect 551910 620509 552230 620593
rect 551910 620273 551952 620509
rect 552188 620273 552230 620509
rect 551910 620241 552230 620273
rect 557840 620829 558160 620861
rect 557840 620593 557882 620829
rect 558118 620593 558160 620829
rect 557840 620509 558160 620593
rect 557840 620273 557882 620509
rect 558118 620273 558160 620509
rect 557840 620241 558160 620273
rect 563771 620829 564091 620861
rect 563771 620593 563813 620829
rect 564049 620593 564091 620829
rect 563771 620509 564091 620593
rect 563771 620273 563813 620509
rect 564049 620273 564091 620509
rect 563771 620241 564091 620273
rect 573494 620829 574114 647273
rect 573494 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 574114 620829
rect 573494 620509 574114 620593
rect 573494 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 574114 620509
rect 22874 617454 23194 617486
rect 22874 617218 22916 617454
rect 23152 617218 23194 617454
rect 22874 617134 23194 617218
rect 22874 616898 22916 617134
rect 23152 616898 23194 617134
rect 22874 616866 23194 616898
rect 28805 617454 29125 617486
rect 28805 617218 28847 617454
rect 29083 617218 29125 617454
rect 28805 617134 29125 617218
rect 28805 616898 28847 617134
rect 29083 616898 29125 617134
rect 28805 616866 29125 616898
rect 50874 617454 51194 617486
rect 50874 617218 50916 617454
rect 51152 617218 51194 617454
rect 50874 617134 51194 617218
rect 50874 616898 50916 617134
rect 51152 616898 51194 617134
rect 50874 616866 51194 616898
rect 56805 617454 57125 617486
rect 56805 617218 56847 617454
rect 57083 617218 57125 617454
rect 56805 617134 57125 617218
rect 56805 616898 56847 617134
rect 57083 616898 57125 617134
rect 56805 616866 57125 616898
rect 78874 617454 79194 617486
rect 78874 617218 78916 617454
rect 79152 617218 79194 617454
rect 78874 617134 79194 617218
rect 78874 616898 78916 617134
rect 79152 616898 79194 617134
rect 78874 616866 79194 616898
rect 84805 617454 85125 617486
rect 84805 617218 84847 617454
rect 85083 617218 85125 617454
rect 84805 617134 85125 617218
rect 84805 616898 84847 617134
rect 85083 616898 85125 617134
rect 84805 616866 85125 616898
rect 106874 617454 107194 617486
rect 106874 617218 106916 617454
rect 107152 617218 107194 617454
rect 106874 617134 107194 617218
rect 106874 616898 106916 617134
rect 107152 616898 107194 617134
rect 106874 616866 107194 616898
rect 112805 617454 113125 617486
rect 112805 617218 112847 617454
rect 113083 617218 113125 617454
rect 112805 617134 113125 617218
rect 112805 616898 112847 617134
rect 113083 616898 113125 617134
rect 112805 616866 113125 616898
rect 134874 617454 135194 617486
rect 134874 617218 134916 617454
rect 135152 617218 135194 617454
rect 134874 617134 135194 617218
rect 134874 616898 134916 617134
rect 135152 616898 135194 617134
rect 134874 616866 135194 616898
rect 140805 617454 141125 617486
rect 140805 617218 140847 617454
rect 141083 617218 141125 617454
rect 140805 617134 141125 617218
rect 140805 616898 140847 617134
rect 141083 616898 141125 617134
rect 140805 616866 141125 616898
rect 162874 617454 163194 617486
rect 162874 617218 162916 617454
rect 163152 617218 163194 617454
rect 162874 617134 163194 617218
rect 162874 616898 162916 617134
rect 163152 616898 163194 617134
rect 162874 616866 163194 616898
rect 168805 617454 169125 617486
rect 168805 617218 168847 617454
rect 169083 617218 169125 617454
rect 168805 617134 169125 617218
rect 168805 616898 168847 617134
rect 169083 616898 169125 617134
rect 168805 616866 169125 616898
rect 190874 617454 191194 617486
rect 190874 617218 190916 617454
rect 191152 617218 191194 617454
rect 190874 617134 191194 617218
rect 190874 616898 190916 617134
rect 191152 616898 191194 617134
rect 190874 616866 191194 616898
rect 196805 617454 197125 617486
rect 196805 617218 196847 617454
rect 197083 617218 197125 617454
rect 196805 617134 197125 617218
rect 196805 616898 196847 617134
rect 197083 616898 197125 617134
rect 196805 616866 197125 616898
rect 218874 617454 219194 617486
rect 218874 617218 218916 617454
rect 219152 617218 219194 617454
rect 218874 617134 219194 617218
rect 218874 616898 218916 617134
rect 219152 616898 219194 617134
rect 218874 616866 219194 616898
rect 224805 617454 225125 617486
rect 224805 617218 224847 617454
rect 225083 617218 225125 617454
rect 224805 617134 225125 617218
rect 224805 616898 224847 617134
rect 225083 616898 225125 617134
rect 224805 616866 225125 616898
rect 246874 617454 247194 617486
rect 246874 617218 246916 617454
rect 247152 617218 247194 617454
rect 246874 617134 247194 617218
rect 246874 616898 246916 617134
rect 247152 616898 247194 617134
rect 246874 616866 247194 616898
rect 252805 617454 253125 617486
rect 252805 617218 252847 617454
rect 253083 617218 253125 617454
rect 252805 617134 253125 617218
rect 252805 616898 252847 617134
rect 253083 616898 253125 617134
rect 252805 616866 253125 616898
rect 274874 617454 275194 617486
rect 274874 617218 274916 617454
rect 275152 617218 275194 617454
rect 274874 617134 275194 617218
rect 274874 616898 274916 617134
rect 275152 616898 275194 617134
rect 274874 616866 275194 616898
rect 280805 617454 281125 617486
rect 280805 617218 280847 617454
rect 281083 617218 281125 617454
rect 280805 617134 281125 617218
rect 280805 616898 280847 617134
rect 281083 616898 281125 617134
rect 280805 616866 281125 616898
rect 302874 617454 303194 617486
rect 302874 617218 302916 617454
rect 303152 617218 303194 617454
rect 302874 617134 303194 617218
rect 302874 616898 302916 617134
rect 303152 616898 303194 617134
rect 302874 616866 303194 616898
rect 308805 617454 309125 617486
rect 308805 617218 308847 617454
rect 309083 617218 309125 617454
rect 308805 617134 309125 617218
rect 308805 616898 308847 617134
rect 309083 616898 309125 617134
rect 308805 616866 309125 616898
rect 330874 617454 331194 617486
rect 330874 617218 330916 617454
rect 331152 617218 331194 617454
rect 330874 617134 331194 617218
rect 330874 616898 330916 617134
rect 331152 616898 331194 617134
rect 330874 616866 331194 616898
rect 336805 617454 337125 617486
rect 336805 617218 336847 617454
rect 337083 617218 337125 617454
rect 336805 617134 337125 617218
rect 336805 616898 336847 617134
rect 337083 616898 337125 617134
rect 336805 616866 337125 616898
rect 358874 617454 359194 617486
rect 358874 617218 358916 617454
rect 359152 617218 359194 617454
rect 358874 617134 359194 617218
rect 358874 616898 358916 617134
rect 359152 616898 359194 617134
rect 358874 616866 359194 616898
rect 364805 617454 365125 617486
rect 364805 617218 364847 617454
rect 365083 617218 365125 617454
rect 364805 617134 365125 617218
rect 364805 616898 364847 617134
rect 365083 616898 365125 617134
rect 364805 616866 365125 616898
rect 386874 617454 387194 617486
rect 386874 617218 386916 617454
rect 387152 617218 387194 617454
rect 386874 617134 387194 617218
rect 386874 616898 386916 617134
rect 387152 616898 387194 617134
rect 386874 616866 387194 616898
rect 392805 617454 393125 617486
rect 392805 617218 392847 617454
rect 393083 617218 393125 617454
rect 392805 617134 393125 617218
rect 392805 616898 392847 617134
rect 393083 616898 393125 617134
rect 392805 616866 393125 616898
rect 414874 617454 415194 617486
rect 414874 617218 414916 617454
rect 415152 617218 415194 617454
rect 414874 617134 415194 617218
rect 414874 616898 414916 617134
rect 415152 616898 415194 617134
rect 414874 616866 415194 616898
rect 420805 617454 421125 617486
rect 420805 617218 420847 617454
rect 421083 617218 421125 617454
rect 420805 617134 421125 617218
rect 420805 616898 420847 617134
rect 421083 616898 421125 617134
rect 420805 616866 421125 616898
rect 442874 617454 443194 617486
rect 442874 617218 442916 617454
rect 443152 617218 443194 617454
rect 442874 617134 443194 617218
rect 442874 616898 442916 617134
rect 443152 616898 443194 617134
rect 442874 616866 443194 616898
rect 448805 617454 449125 617486
rect 448805 617218 448847 617454
rect 449083 617218 449125 617454
rect 448805 617134 449125 617218
rect 448805 616898 448847 617134
rect 449083 616898 449125 617134
rect 448805 616866 449125 616898
rect 470874 617454 471194 617486
rect 470874 617218 470916 617454
rect 471152 617218 471194 617454
rect 470874 617134 471194 617218
rect 470874 616898 470916 617134
rect 471152 616898 471194 617134
rect 470874 616866 471194 616898
rect 476805 617454 477125 617486
rect 476805 617218 476847 617454
rect 477083 617218 477125 617454
rect 476805 617134 477125 617218
rect 476805 616898 476847 617134
rect 477083 616898 477125 617134
rect 476805 616866 477125 616898
rect 498874 617454 499194 617486
rect 498874 617218 498916 617454
rect 499152 617218 499194 617454
rect 498874 617134 499194 617218
rect 498874 616898 498916 617134
rect 499152 616898 499194 617134
rect 498874 616866 499194 616898
rect 504805 617454 505125 617486
rect 504805 617218 504847 617454
rect 505083 617218 505125 617454
rect 504805 617134 505125 617218
rect 504805 616898 504847 617134
rect 505083 616898 505125 617134
rect 504805 616866 505125 616898
rect 526874 617454 527194 617486
rect 526874 617218 526916 617454
rect 527152 617218 527194 617454
rect 526874 617134 527194 617218
rect 526874 616898 526916 617134
rect 527152 616898 527194 617134
rect 526874 616866 527194 616898
rect 532805 617454 533125 617486
rect 532805 617218 532847 617454
rect 533083 617218 533125 617454
rect 532805 617134 533125 617218
rect 532805 616898 532847 617134
rect 533083 616898 533125 617134
rect 532805 616866 533125 616898
rect 554874 617454 555194 617486
rect 554874 617218 554916 617454
rect 555152 617218 555194 617454
rect 554874 617134 555194 617218
rect 554874 616898 554916 617134
rect 555152 616898 555194 617134
rect 554874 616866 555194 616898
rect 560805 617454 561125 617486
rect 560805 617218 560847 617454
rect 561083 617218 561125 617454
rect 560805 617134 561125 617218
rect 560805 616898 560847 617134
rect 561083 616898 561125 617134
rect 560805 616866 561125 616898
rect -2006 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 -1386 593829
rect -2006 593509 -1386 593593
rect -2006 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 -1386 593509
rect -2006 566829 -1386 593273
rect 19910 593829 20230 593861
rect 19910 593593 19952 593829
rect 20188 593593 20230 593829
rect 19910 593509 20230 593593
rect 19910 593273 19952 593509
rect 20188 593273 20230 593509
rect 19910 593241 20230 593273
rect 25840 593829 26160 593861
rect 25840 593593 25882 593829
rect 26118 593593 26160 593829
rect 25840 593509 26160 593593
rect 25840 593273 25882 593509
rect 26118 593273 26160 593509
rect 25840 593241 26160 593273
rect 31771 593829 32091 593861
rect 31771 593593 31813 593829
rect 32049 593593 32091 593829
rect 31771 593509 32091 593593
rect 31771 593273 31813 593509
rect 32049 593273 32091 593509
rect 31771 593241 32091 593273
rect 47910 593829 48230 593861
rect 47910 593593 47952 593829
rect 48188 593593 48230 593829
rect 47910 593509 48230 593593
rect 47910 593273 47952 593509
rect 48188 593273 48230 593509
rect 47910 593241 48230 593273
rect 53840 593829 54160 593861
rect 53840 593593 53882 593829
rect 54118 593593 54160 593829
rect 53840 593509 54160 593593
rect 53840 593273 53882 593509
rect 54118 593273 54160 593509
rect 53840 593241 54160 593273
rect 59771 593829 60091 593861
rect 59771 593593 59813 593829
rect 60049 593593 60091 593829
rect 59771 593509 60091 593593
rect 59771 593273 59813 593509
rect 60049 593273 60091 593509
rect 59771 593241 60091 593273
rect 75910 593829 76230 593861
rect 75910 593593 75952 593829
rect 76188 593593 76230 593829
rect 75910 593509 76230 593593
rect 75910 593273 75952 593509
rect 76188 593273 76230 593509
rect 75910 593241 76230 593273
rect 81840 593829 82160 593861
rect 81840 593593 81882 593829
rect 82118 593593 82160 593829
rect 81840 593509 82160 593593
rect 81840 593273 81882 593509
rect 82118 593273 82160 593509
rect 81840 593241 82160 593273
rect 87771 593829 88091 593861
rect 87771 593593 87813 593829
rect 88049 593593 88091 593829
rect 87771 593509 88091 593593
rect 87771 593273 87813 593509
rect 88049 593273 88091 593509
rect 87771 593241 88091 593273
rect 103910 593829 104230 593861
rect 103910 593593 103952 593829
rect 104188 593593 104230 593829
rect 103910 593509 104230 593593
rect 103910 593273 103952 593509
rect 104188 593273 104230 593509
rect 103910 593241 104230 593273
rect 109840 593829 110160 593861
rect 109840 593593 109882 593829
rect 110118 593593 110160 593829
rect 109840 593509 110160 593593
rect 109840 593273 109882 593509
rect 110118 593273 110160 593509
rect 109840 593241 110160 593273
rect 115771 593829 116091 593861
rect 115771 593593 115813 593829
rect 116049 593593 116091 593829
rect 115771 593509 116091 593593
rect 115771 593273 115813 593509
rect 116049 593273 116091 593509
rect 115771 593241 116091 593273
rect 131910 593829 132230 593861
rect 131910 593593 131952 593829
rect 132188 593593 132230 593829
rect 131910 593509 132230 593593
rect 131910 593273 131952 593509
rect 132188 593273 132230 593509
rect 131910 593241 132230 593273
rect 137840 593829 138160 593861
rect 137840 593593 137882 593829
rect 138118 593593 138160 593829
rect 137840 593509 138160 593593
rect 137840 593273 137882 593509
rect 138118 593273 138160 593509
rect 137840 593241 138160 593273
rect 143771 593829 144091 593861
rect 143771 593593 143813 593829
rect 144049 593593 144091 593829
rect 143771 593509 144091 593593
rect 143771 593273 143813 593509
rect 144049 593273 144091 593509
rect 143771 593241 144091 593273
rect 159910 593829 160230 593861
rect 159910 593593 159952 593829
rect 160188 593593 160230 593829
rect 159910 593509 160230 593593
rect 159910 593273 159952 593509
rect 160188 593273 160230 593509
rect 159910 593241 160230 593273
rect 165840 593829 166160 593861
rect 165840 593593 165882 593829
rect 166118 593593 166160 593829
rect 165840 593509 166160 593593
rect 165840 593273 165882 593509
rect 166118 593273 166160 593509
rect 165840 593241 166160 593273
rect 171771 593829 172091 593861
rect 171771 593593 171813 593829
rect 172049 593593 172091 593829
rect 171771 593509 172091 593593
rect 171771 593273 171813 593509
rect 172049 593273 172091 593509
rect 171771 593241 172091 593273
rect 187910 593829 188230 593861
rect 187910 593593 187952 593829
rect 188188 593593 188230 593829
rect 187910 593509 188230 593593
rect 187910 593273 187952 593509
rect 188188 593273 188230 593509
rect 187910 593241 188230 593273
rect 193840 593829 194160 593861
rect 193840 593593 193882 593829
rect 194118 593593 194160 593829
rect 193840 593509 194160 593593
rect 193840 593273 193882 593509
rect 194118 593273 194160 593509
rect 193840 593241 194160 593273
rect 199771 593829 200091 593861
rect 199771 593593 199813 593829
rect 200049 593593 200091 593829
rect 199771 593509 200091 593593
rect 199771 593273 199813 593509
rect 200049 593273 200091 593509
rect 199771 593241 200091 593273
rect 215910 593829 216230 593861
rect 215910 593593 215952 593829
rect 216188 593593 216230 593829
rect 215910 593509 216230 593593
rect 215910 593273 215952 593509
rect 216188 593273 216230 593509
rect 215910 593241 216230 593273
rect 221840 593829 222160 593861
rect 221840 593593 221882 593829
rect 222118 593593 222160 593829
rect 221840 593509 222160 593593
rect 221840 593273 221882 593509
rect 222118 593273 222160 593509
rect 221840 593241 222160 593273
rect 227771 593829 228091 593861
rect 227771 593593 227813 593829
rect 228049 593593 228091 593829
rect 227771 593509 228091 593593
rect 227771 593273 227813 593509
rect 228049 593273 228091 593509
rect 227771 593241 228091 593273
rect 243910 593829 244230 593861
rect 243910 593593 243952 593829
rect 244188 593593 244230 593829
rect 243910 593509 244230 593593
rect 243910 593273 243952 593509
rect 244188 593273 244230 593509
rect 243910 593241 244230 593273
rect 249840 593829 250160 593861
rect 249840 593593 249882 593829
rect 250118 593593 250160 593829
rect 249840 593509 250160 593593
rect 249840 593273 249882 593509
rect 250118 593273 250160 593509
rect 249840 593241 250160 593273
rect 255771 593829 256091 593861
rect 255771 593593 255813 593829
rect 256049 593593 256091 593829
rect 255771 593509 256091 593593
rect 255771 593273 255813 593509
rect 256049 593273 256091 593509
rect 255771 593241 256091 593273
rect 271910 593829 272230 593861
rect 271910 593593 271952 593829
rect 272188 593593 272230 593829
rect 271910 593509 272230 593593
rect 271910 593273 271952 593509
rect 272188 593273 272230 593509
rect 271910 593241 272230 593273
rect 277840 593829 278160 593861
rect 277840 593593 277882 593829
rect 278118 593593 278160 593829
rect 277840 593509 278160 593593
rect 277840 593273 277882 593509
rect 278118 593273 278160 593509
rect 277840 593241 278160 593273
rect 283771 593829 284091 593861
rect 283771 593593 283813 593829
rect 284049 593593 284091 593829
rect 283771 593509 284091 593593
rect 283771 593273 283813 593509
rect 284049 593273 284091 593509
rect 283771 593241 284091 593273
rect 299910 593829 300230 593861
rect 299910 593593 299952 593829
rect 300188 593593 300230 593829
rect 299910 593509 300230 593593
rect 299910 593273 299952 593509
rect 300188 593273 300230 593509
rect 299910 593241 300230 593273
rect 305840 593829 306160 593861
rect 305840 593593 305882 593829
rect 306118 593593 306160 593829
rect 305840 593509 306160 593593
rect 305840 593273 305882 593509
rect 306118 593273 306160 593509
rect 305840 593241 306160 593273
rect 311771 593829 312091 593861
rect 311771 593593 311813 593829
rect 312049 593593 312091 593829
rect 311771 593509 312091 593593
rect 311771 593273 311813 593509
rect 312049 593273 312091 593509
rect 311771 593241 312091 593273
rect 327910 593829 328230 593861
rect 327910 593593 327952 593829
rect 328188 593593 328230 593829
rect 327910 593509 328230 593593
rect 327910 593273 327952 593509
rect 328188 593273 328230 593509
rect 327910 593241 328230 593273
rect 333840 593829 334160 593861
rect 333840 593593 333882 593829
rect 334118 593593 334160 593829
rect 333840 593509 334160 593593
rect 333840 593273 333882 593509
rect 334118 593273 334160 593509
rect 333840 593241 334160 593273
rect 339771 593829 340091 593861
rect 339771 593593 339813 593829
rect 340049 593593 340091 593829
rect 339771 593509 340091 593593
rect 339771 593273 339813 593509
rect 340049 593273 340091 593509
rect 339771 593241 340091 593273
rect 355910 593829 356230 593861
rect 355910 593593 355952 593829
rect 356188 593593 356230 593829
rect 355910 593509 356230 593593
rect 355910 593273 355952 593509
rect 356188 593273 356230 593509
rect 355910 593241 356230 593273
rect 361840 593829 362160 593861
rect 361840 593593 361882 593829
rect 362118 593593 362160 593829
rect 361840 593509 362160 593593
rect 361840 593273 361882 593509
rect 362118 593273 362160 593509
rect 361840 593241 362160 593273
rect 367771 593829 368091 593861
rect 367771 593593 367813 593829
rect 368049 593593 368091 593829
rect 367771 593509 368091 593593
rect 367771 593273 367813 593509
rect 368049 593273 368091 593509
rect 367771 593241 368091 593273
rect 383910 593829 384230 593861
rect 383910 593593 383952 593829
rect 384188 593593 384230 593829
rect 383910 593509 384230 593593
rect 383910 593273 383952 593509
rect 384188 593273 384230 593509
rect 383910 593241 384230 593273
rect 389840 593829 390160 593861
rect 389840 593593 389882 593829
rect 390118 593593 390160 593829
rect 389840 593509 390160 593593
rect 389840 593273 389882 593509
rect 390118 593273 390160 593509
rect 389840 593241 390160 593273
rect 395771 593829 396091 593861
rect 395771 593593 395813 593829
rect 396049 593593 396091 593829
rect 395771 593509 396091 593593
rect 395771 593273 395813 593509
rect 396049 593273 396091 593509
rect 395771 593241 396091 593273
rect 411910 593829 412230 593861
rect 411910 593593 411952 593829
rect 412188 593593 412230 593829
rect 411910 593509 412230 593593
rect 411910 593273 411952 593509
rect 412188 593273 412230 593509
rect 411910 593241 412230 593273
rect 417840 593829 418160 593861
rect 417840 593593 417882 593829
rect 418118 593593 418160 593829
rect 417840 593509 418160 593593
rect 417840 593273 417882 593509
rect 418118 593273 418160 593509
rect 417840 593241 418160 593273
rect 423771 593829 424091 593861
rect 423771 593593 423813 593829
rect 424049 593593 424091 593829
rect 423771 593509 424091 593593
rect 423771 593273 423813 593509
rect 424049 593273 424091 593509
rect 423771 593241 424091 593273
rect 439910 593829 440230 593861
rect 439910 593593 439952 593829
rect 440188 593593 440230 593829
rect 439910 593509 440230 593593
rect 439910 593273 439952 593509
rect 440188 593273 440230 593509
rect 439910 593241 440230 593273
rect 445840 593829 446160 593861
rect 445840 593593 445882 593829
rect 446118 593593 446160 593829
rect 445840 593509 446160 593593
rect 445840 593273 445882 593509
rect 446118 593273 446160 593509
rect 445840 593241 446160 593273
rect 451771 593829 452091 593861
rect 451771 593593 451813 593829
rect 452049 593593 452091 593829
rect 451771 593509 452091 593593
rect 451771 593273 451813 593509
rect 452049 593273 452091 593509
rect 451771 593241 452091 593273
rect 467910 593829 468230 593861
rect 467910 593593 467952 593829
rect 468188 593593 468230 593829
rect 467910 593509 468230 593593
rect 467910 593273 467952 593509
rect 468188 593273 468230 593509
rect 467910 593241 468230 593273
rect 473840 593829 474160 593861
rect 473840 593593 473882 593829
rect 474118 593593 474160 593829
rect 473840 593509 474160 593593
rect 473840 593273 473882 593509
rect 474118 593273 474160 593509
rect 473840 593241 474160 593273
rect 479771 593829 480091 593861
rect 479771 593593 479813 593829
rect 480049 593593 480091 593829
rect 479771 593509 480091 593593
rect 479771 593273 479813 593509
rect 480049 593273 480091 593509
rect 479771 593241 480091 593273
rect 495910 593829 496230 593861
rect 495910 593593 495952 593829
rect 496188 593593 496230 593829
rect 495910 593509 496230 593593
rect 495910 593273 495952 593509
rect 496188 593273 496230 593509
rect 495910 593241 496230 593273
rect 501840 593829 502160 593861
rect 501840 593593 501882 593829
rect 502118 593593 502160 593829
rect 501840 593509 502160 593593
rect 501840 593273 501882 593509
rect 502118 593273 502160 593509
rect 501840 593241 502160 593273
rect 507771 593829 508091 593861
rect 507771 593593 507813 593829
rect 508049 593593 508091 593829
rect 507771 593509 508091 593593
rect 507771 593273 507813 593509
rect 508049 593273 508091 593509
rect 507771 593241 508091 593273
rect 523910 593829 524230 593861
rect 523910 593593 523952 593829
rect 524188 593593 524230 593829
rect 523910 593509 524230 593593
rect 523910 593273 523952 593509
rect 524188 593273 524230 593509
rect 523910 593241 524230 593273
rect 529840 593829 530160 593861
rect 529840 593593 529882 593829
rect 530118 593593 530160 593829
rect 529840 593509 530160 593593
rect 529840 593273 529882 593509
rect 530118 593273 530160 593509
rect 529840 593241 530160 593273
rect 535771 593829 536091 593861
rect 535771 593593 535813 593829
rect 536049 593593 536091 593829
rect 535771 593509 536091 593593
rect 535771 593273 535813 593509
rect 536049 593273 536091 593509
rect 535771 593241 536091 593273
rect 551910 593829 552230 593861
rect 551910 593593 551952 593829
rect 552188 593593 552230 593829
rect 551910 593509 552230 593593
rect 551910 593273 551952 593509
rect 552188 593273 552230 593509
rect 551910 593241 552230 593273
rect 557840 593829 558160 593861
rect 557840 593593 557882 593829
rect 558118 593593 558160 593829
rect 557840 593509 558160 593593
rect 557840 593273 557882 593509
rect 558118 593273 558160 593509
rect 557840 593241 558160 593273
rect 563771 593829 564091 593861
rect 563771 593593 563813 593829
rect 564049 593593 564091 593829
rect 563771 593509 564091 593593
rect 563771 593273 563813 593509
rect 564049 593273 564091 593509
rect 563771 593241 564091 593273
rect 573494 593829 574114 620273
rect 573494 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 574114 593829
rect 573494 593509 574114 593593
rect 573494 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 574114 593509
rect 22874 590454 23194 590486
rect 22874 590218 22916 590454
rect 23152 590218 23194 590454
rect 22874 590134 23194 590218
rect 22874 589898 22916 590134
rect 23152 589898 23194 590134
rect 22874 589866 23194 589898
rect 28805 590454 29125 590486
rect 28805 590218 28847 590454
rect 29083 590218 29125 590454
rect 28805 590134 29125 590218
rect 28805 589898 28847 590134
rect 29083 589898 29125 590134
rect 28805 589866 29125 589898
rect 50874 590454 51194 590486
rect 50874 590218 50916 590454
rect 51152 590218 51194 590454
rect 50874 590134 51194 590218
rect 50874 589898 50916 590134
rect 51152 589898 51194 590134
rect 50874 589866 51194 589898
rect 56805 590454 57125 590486
rect 56805 590218 56847 590454
rect 57083 590218 57125 590454
rect 56805 590134 57125 590218
rect 56805 589898 56847 590134
rect 57083 589898 57125 590134
rect 56805 589866 57125 589898
rect 78874 590454 79194 590486
rect 78874 590218 78916 590454
rect 79152 590218 79194 590454
rect 78874 590134 79194 590218
rect 78874 589898 78916 590134
rect 79152 589898 79194 590134
rect 78874 589866 79194 589898
rect 84805 590454 85125 590486
rect 84805 590218 84847 590454
rect 85083 590218 85125 590454
rect 84805 590134 85125 590218
rect 84805 589898 84847 590134
rect 85083 589898 85125 590134
rect 84805 589866 85125 589898
rect 106874 590454 107194 590486
rect 106874 590218 106916 590454
rect 107152 590218 107194 590454
rect 106874 590134 107194 590218
rect 106874 589898 106916 590134
rect 107152 589898 107194 590134
rect 106874 589866 107194 589898
rect 112805 590454 113125 590486
rect 112805 590218 112847 590454
rect 113083 590218 113125 590454
rect 112805 590134 113125 590218
rect 112805 589898 112847 590134
rect 113083 589898 113125 590134
rect 112805 589866 113125 589898
rect 134874 590454 135194 590486
rect 134874 590218 134916 590454
rect 135152 590218 135194 590454
rect 134874 590134 135194 590218
rect 134874 589898 134916 590134
rect 135152 589898 135194 590134
rect 134874 589866 135194 589898
rect 140805 590454 141125 590486
rect 140805 590218 140847 590454
rect 141083 590218 141125 590454
rect 140805 590134 141125 590218
rect 140805 589898 140847 590134
rect 141083 589898 141125 590134
rect 140805 589866 141125 589898
rect 162874 590454 163194 590486
rect 162874 590218 162916 590454
rect 163152 590218 163194 590454
rect 162874 590134 163194 590218
rect 162874 589898 162916 590134
rect 163152 589898 163194 590134
rect 162874 589866 163194 589898
rect 168805 590454 169125 590486
rect 168805 590218 168847 590454
rect 169083 590218 169125 590454
rect 168805 590134 169125 590218
rect 168805 589898 168847 590134
rect 169083 589898 169125 590134
rect 168805 589866 169125 589898
rect 190874 590454 191194 590486
rect 190874 590218 190916 590454
rect 191152 590218 191194 590454
rect 190874 590134 191194 590218
rect 190874 589898 190916 590134
rect 191152 589898 191194 590134
rect 190874 589866 191194 589898
rect 196805 590454 197125 590486
rect 196805 590218 196847 590454
rect 197083 590218 197125 590454
rect 196805 590134 197125 590218
rect 196805 589898 196847 590134
rect 197083 589898 197125 590134
rect 196805 589866 197125 589898
rect 218874 590454 219194 590486
rect 218874 590218 218916 590454
rect 219152 590218 219194 590454
rect 218874 590134 219194 590218
rect 218874 589898 218916 590134
rect 219152 589898 219194 590134
rect 218874 589866 219194 589898
rect 224805 590454 225125 590486
rect 224805 590218 224847 590454
rect 225083 590218 225125 590454
rect 224805 590134 225125 590218
rect 224805 589898 224847 590134
rect 225083 589898 225125 590134
rect 224805 589866 225125 589898
rect 246874 590454 247194 590486
rect 246874 590218 246916 590454
rect 247152 590218 247194 590454
rect 246874 590134 247194 590218
rect 246874 589898 246916 590134
rect 247152 589898 247194 590134
rect 246874 589866 247194 589898
rect 252805 590454 253125 590486
rect 252805 590218 252847 590454
rect 253083 590218 253125 590454
rect 252805 590134 253125 590218
rect 252805 589898 252847 590134
rect 253083 589898 253125 590134
rect 252805 589866 253125 589898
rect 274874 590454 275194 590486
rect 274874 590218 274916 590454
rect 275152 590218 275194 590454
rect 274874 590134 275194 590218
rect 274874 589898 274916 590134
rect 275152 589898 275194 590134
rect 274874 589866 275194 589898
rect 280805 590454 281125 590486
rect 280805 590218 280847 590454
rect 281083 590218 281125 590454
rect 280805 590134 281125 590218
rect 280805 589898 280847 590134
rect 281083 589898 281125 590134
rect 280805 589866 281125 589898
rect 302874 590454 303194 590486
rect 302874 590218 302916 590454
rect 303152 590218 303194 590454
rect 302874 590134 303194 590218
rect 302874 589898 302916 590134
rect 303152 589898 303194 590134
rect 302874 589866 303194 589898
rect 308805 590454 309125 590486
rect 308805 590218 308847 590454
rect 309083 590218 309125 590454
rect 308805 590134 309125 590218
rect 308805 589898 308847 590134
rect 309083 589898 309125 590134
rect 308805 589866 309125 589898
rect 330874 590454 331194 590486
rect 330874 590218 330916 590454
rect 331152 590218 331194 590454
rect 330874 590134 331194 590218
rect 330874 589898 330916 590134
rect 331152 589898 331194 590134
rect 330874 589866 331194 589898
rect 336805 590454 337125 590486
rect 336805 590218 336847 590454
rect 337083 590218 337125 590454
rect 336805 590134 337125 590218
rect 336805 589898 336847 590134
rect 337083 589898 337125 590134
rect 336805 589866 337125 589898
rect 358874 590454 359194 590486
rect 358874 590218 358916 590454
rect 359152 590218 359194 590454
rect 358874 590134 359194 590218
rect 358874 589898 358916 590134
rect 359152 589898 359194 590134
rect 358874 589866 359194 589898
rect 364805 590454 365125 590486
rect 364805 590218 364847 590454
rect 365083 590218 365125 590454
rect 364805 590134 365125 590218
rect 364805 589898 364847 590134
rect 365083 589898 365125 590134
rect 364805 589866 365125 589898
rect 386874 590454 387194 590486
rect 386874 590218 386916 590454
rect 387152 590218 387194 590454
rect 386874 590134 387194 590218
rect 386874 589898 386916 590134
rect 387152 589898 387194 590134
rect 386874 589866 387194 589898
rect 392805 590454 393125 590486
rect 392805 590218 392847 590454
rect 393083 590218 393125 590454
rect 392805 590134 393125 590218
rect 392805 589898 392847 590134
rect 393083 589898 393125 590134
rect 392805 589866 393125 589898
rect 414874 590454 415194 590486
rect 414874 590218 414916 590454
rect 415152 590218 415194 590454
rect 414874 590134 415194 590218
rect 414874 589898 414916 590134
rect 415152 589898 415194 590134
rect 414874 589866 415194 589898
rect 420805 590454 421125 590486
rect 420805 590218 420847 590454
rect 421083 590218 421125 590454
rect 420805 590134 421125 590218
rect 420805 589898 420847 590134
rect 421083 589898 421125 590134
rect 420805 589866 421125 589898
rect 442874 590454 443194 590486
rect 442874 590218 442916 590454
rect 443152 590218 443194 590454
rect 442874 590134 443194 590218
rect 442874 589898 442916 590134
rect 443152 589898 443194 590134
rect 442874 589866 443194 589898
rect 448805 590454 449125 590486
rect 448805 590218 448847 590454
rect 449083 590218 449125 590454
rect 448805 590134 449125 590218
rect 448805 589898 448847 590134
rect 449083 589898 449125 590134
rect 448805 589866 449125 589898
rect 470874 590454 471194 590486
rect 470874 590218 470916 590454
rect 471152 590218 471194 590454
rect 470874 590134 471194 590218
rect 470874 589898 470916 590134
rect 471152 589898 471194 590134
rect 470874 589866 471194 589898
rect 476805 590454 477125 590486
rect 476805 590218 476847 590454
rect 477083 590218 477125 590454
rect 476805 590134 477125 590218
rect 476805 589898 476847 590134
rect 477083 589898 477125 590134
rect 476805 589866 477125 589898
rect 498874 590454 499194 590486
rect 498874 590218 498916 590454
rect 499152 590218 499194 590454
rect 498874 590134 499194 590218
rect 498874 589898 498916 590134
rect 499152 589898 499194 590134
rect 498874 589866 499194 589898
rect 504805 590454 505125 590486
rect 504805 590218 504847 590454
rect 505083 590218 505125 590454
rect 504805 590134 505125 590218
rect 504805 589898 504847 590134
rect 505083 589898 505125 590134
rect 504805 589866 505125 589898
rect 526874 590454 527194 590486
rect 526874 590218 526916 590454
rect 527152 590218 527194 590454
rect 526874 590134 527194 590218
rect 526874 589898 526916 590134
rect 527152 589898 527194 590134
rect 526874 589866 527194 589898
rect 532805 590454 533125 590486
rect 532805 590218 532847 590454
rect 533083 590218 533125 590454
rect 532805 590134 533125 590218
rect 532805 589898 532847 590134
rect 533083 589898 533125 590134
rect 532805 589866 533125 589898
rect 554874 590454 555194 590486
rect 554874 590218 554916 590454
rect 555152 590218 555194 590454
rect 554874 590134 555194 590218
rect 554874 589898 554916 590134
rect 555152 589898 555194 590134
rect 554874 589866 555194 589898
rect 560805 590454 561125 590486
rect 560805 590218 560847 590454
rect 561083 590218 561125 590454
rect 560805 590134 561125 590218
rect 560805 589898 560847 590134
rect 561083 589898 561125 590134
rect 560805 589866 561125 589898
rect -2006 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 -1386 566829
rect -2006 566509 -1386 566593
rect -2006 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 -1386 566509
rect -2006 539829 -1386 566273
rect 19910 566829 20230 566861
rect 19910 566593 19952 566829
rect 20188 566593 20230 566829
rect 19910 566509 20230 566593
rect 19910 566273 19952 566509
rect 20188 566273 20230 566509
rect 19910 566241 20230 566273
rect 25840 566829 26160 566861
rect 25840 566593 25882 566829
rect 26118 566593 26160 566829
rect 25840 566509 26160 566593
rect 25840 566273 25882 566509
rect 26118 566273 26160 566509
rect 25840 566241 26160 566273
rect 31771 566829 32091 566861
rect 31771 566593 31813 566829
rect 32049 566593 32091 566829
rect 31771 566509 32091 566593
rect 31771 566273 31813 566509
rect 32049 566273 32091 566509
rect 31771 566241 32091 566273
rect 47910 566829 48230 566861
rect 47910 566593 47952 566829
rect 48188 566593 48230 566829
rect 47910 566509 48230 566593
rect 47910 566273 47952 566509
rect 48188 566273 48230 566509
rect 47910 566241 48230 566273
rect 53840 566829 54160 566861
rect 53840 566593 53882 566829
rect 54118 566593 54160 566829
rect 53840 566509 54160 566593
rect 53840 566273 53882 566509
rect 54118 566273 54160 566509
rect 53840 566241 54160 566273
rect 59771 566829 60091 566861
rect 59771 566593 59813 566829
rect 60049 566593 60091 566829
rect 59771 566509 60091 566593
rect 59771 566273 59813 566509
rect 60049 566273 60091 566509
rect 59771 566241 60091 566273
rect 75910 566829 76230 566861
rect 75910 566593 75952 566829
rect 76188 566593 76230 566829
rect 75910 566509 76230 566593
rect 75910 566273 75952 566509
rect 76188 566273 76230 566509
rect 75910 566241 76230 566273
rect 81840 566829 82160 566861
rect 81840 566593 81882 566829
rect 82118 566593 82160 566829
rect 81840 566509 82160 566593
rect 81840 566273 81882 566509
rect 82118 566273 82160 566509
rect 81840 566241 82160 566273
rect 87771 566829 88091 566861
rect 87771 566593 87813 566829
rect 88049 566593 88091 566829
rect 87771 566509 88091 566593
rect 87771 566273 87813 566509
rect 88049 566273 88091 566509
rect 87771 566241 88091 566273
rect 103910 566829 104230 566861
rect 103910 566593 103952 566829
rect 104188 566593 104230 566829
rect 103910 566509 104230 566593
rect 103910 566273 103952 566509
rect 104188 566273 104230 566509
rect 103910 566241 104230 566273
rect 109840 566829 110160 566861
rect 109840 566593 109882 566829
rect 110118 566593 110160 566829
rect 109840 566509 110160 566593
rect 109840 566273 109882 566509
rect 110118 566273 110160 566509
rect 109840 566241 110160 566273
rect 115771 566829 116091 566861
rect 115771 566593 115813 566829
rect 116049 566593 116091 566829
rect 115771 566509 116091 566593
rect 115771 566273 115813 566509
rect 116049 566273 116091 566509
rect 115771 566241 116091 566273
rect 131910 566829 132230 566861
rect 131910 566593 131952 566829
rect 132188 566593 132230 566829
rect 131910 566509 132230 566593
rect 131910 566273 131952 566509
rect 132188 566273 132230 566509
rect 131910 566241 132230 566273
rect 137840 566829 138160 566861
rect 137840 566593 137882 566829
rect 138118 566593 138160 566829
rect 137840 566509 138160 566593
rect 137840 566273 137882 566509
rect 138118 566273 138160 566509
rect 137840 566241 138160 566273
rect 143771 566829 144091 566861
rect 143771 566593 143813 566829
rect 144049 566593 144091 566829
rect 143771 566509 144091 566593
rect 143771 566273 143813 566509
rect 144049 566273 144091 566509
rect 143771 566241 144091 566273
rect 159910 566829 160230 566861
rect 159910 566593 159952 566829
rect 160188 566593 160230 566829
rect 159910 566509 160230 566593
rect 159910 566273 159952 566509
rect 160188 566273 160230 566509
rect 159910 566241 160230 566273
rect 165840 566829 166160 566861
rect 165840 566593 165882 566829
rect 166118 566593 166160 566829
rect 165840 566509 166160 566593
rect 165840 566273 165882 566509
rect 166118 566273 166160 566509
rect 165840 566241 166160 566273
rect 171771 566829 172091 566861
rect 171771 566593 171813 566829
rect 172049 566593 172091 566829
rect 171771 566509 172091 566593
rect 171771 566273 171813 566509
rect 172049 566273 172091 566509
rect 171771 566241 172091 566273
rect 187910 566829 188230 566861
rect 187910 566593 187952 566829
rect 188188 566593 188230 566829
rect 187910 566509 188230 566593
rect 187910 566273 187952 566509
rect 188188 566273 188230 566509
rect 187910 566241 188230 566273
rect 193840 566829 194160 566861
rect 193840 566593 193882 566829
rect 194118 566593 194160 566829
rect 193840 566509 194160 566593
rect 193840 566273 193882 566509
rect 194118 566273 194160 566509
rect 193840 566241 194160 566273
rect 199771 566829 200091 566861
rect 199771 566593 199813 566829
rect 200049 566593 200091 566829
rect 199771 566509 200091 566593
rect 199771 566273 199813 566509
rect 200049 566273 200091 566509
rect 199771 566241 200091 566273
rect 215910 566829 216230 566861
rect 215910 566593 215952 566829
rect 216188 566593 216230 566829
rect 215910 566509 216230 566593
rect 215910 566273 215952 566509
rect 216188 566273 216230 566509
rect 215910 566241 216230 566273
rect 221840 566829 222160 566861
rect 221840 566593 221882 566829
rect 222118 566593 222160 566829
rect 221840 566509 222160 566593
rect 221840 566273 221882 566509
rect 222118 566273 222160 566509
rect 221840 566241 222160 566273
rect 227771 566829 228091 566861
rect 227771 566593 227813 566829
rect 228049 566593 228091 566829
rect 227771 566509 228091 566593
rect 227771 566273 227813 566509
rect 228049 566273 228091 566509
rect 227771 566241 228091 566273
rect 243910 566829 244230 566861
rect 243910 566593 243952 566829
rect 244188 566593 244230 566829
rect 243910 566509 244230 566593
rect 243910 566273 243952 566509
rect 244188 566273 244230 566509
rect 243910 566241 244230 566273
rect 249840 566829 250160 566861
rect 249840 566593 249882 566829
rect 250118 566593 250160 566829
rect 249840 566509 250160 566593
rect 249840 566273 249882 566509
rect 250118 566273 250160 566509
rect 249840 566241 250160 566273
rect 255771 566829 256091 566861
rect 255771 566593 255813 566829
rect 256049 566593 256091 566829
rect 255771 566509 256091 566593
rect 255771 566273 255813 566509
rect 256049 566273 256091 566509
rect 255771 566241 256091 566273
rect 271910 566829 272230 566861
rect 271910 566593 271952 566829
rect 272188 566593 272230 566829
rect 271910 566509 272230 566593
rect 271910 566273 271952 566509
rect 272188 566273 272230 566509
rect 271910 566241 272230 566273
rect 277840 566829 278160 566861
rect 277840 566593 277882 566829
rect 278118 566593 278160 566829
rect 277840 566509 278160 566593
rect 277840 566273 277882 566509
rect 278118 566273 278160 566509
rect 277840 566241 278160 566273
rect 283771 566829 284091 566861
rect 283771 566593 283813 566829
rect 284049 566593 284091 566829
rect 283771 566509 284091 566593
rect 283771 566273 283813 566509
rect 284049 566273 284091 566509
rect 283771 566241 284091 566273
rect 299910 566829 300230 566861
rect 299910 566593 299952 566829
rect 300188 566593 300230 566829
rect 299910 566509 300230 566593
rect 299910 566273 299952 566509
rect 300188 566273 300230 566509
rect 299910 566241 300230 566273
rect 305840 566829 306160 566861
rect 305840 566593 305882 566829
rect 306118 566593 306160 566829
rect 305840 566509 306160 566593
rect 305840 566273 305882 566509
rect 306118 566273 306160 566509
rect 305840 566241 306160 566273
rect 311771 566829 312091 566861
rect 311771 566593 311813 566829
rect 312049 566593 312091 566829
rect 311771 566509 312091 566593
rect 311771 566273 311813 566509
rect 312049 566273 312091 566509
rect 311771 566241 312091 566273
rect 327910 566829 328230 566861
rect 327910 566593 327952 566829
rect 328188 566593 328230 566829
rect 327910 566509 328230 566593
rect 327910 566273 327952 566509
rect 328188 566273 328230 566509
rect 327910 566241 328230 566273
rect 333840 566829 334160 566861
rect 333840 566593 333882 566829
rect 334118 566593 334160 566829
rect 333840 566509 334160 566593
rect 333840 566273 333882 566509
rect 334118 566273 334160 566509
rect 333840 566241 334160 566273
rect 339771 566829 340091 566861
rect 339771 566593 339813 566829
rect 340049 566593 340091 566829
rect 339771 566509 340091 566593
rect 339771 566273 339813 566509
rect 340049 566273 340091 566509
rect 339771 566241 340091 566273
rect 355910 566829 356230 566861
rect 355910 566593 355952 566829
rect 356188 566593 356230 566829
rect 355910 566509 356230 566593
rect 355910 566273 355952 566509
rect 356188 566273 356230 566509
rect 355910 566241 356230 566273
rect 361840 566829 362160 566861
rect 361840 566593 361882 566829
rect 362118 566593 362160 566829
rect 361840 566509 362160 566593
rect 361840 566273 361882 566509
rect 362118 566273 362160 566509
rect 361840 566241 362160 566273
rect 367771 566829 368091 566861
rect 367771 566593 367813 566829
rect 368049 566593 368091 566829
rect 367771 566509 368091 566593
rect 367771 566273 367813 566509
rect 368049 566273 368091 566509
rect 367771 566241 368091 566273
rect 383910 566829 384230 566861
rect 383910 566593 383952 566829
rect 384188 566593 384230 566829
rect 383910 566509 384230 566593
rect 383910 566273 383952 566509
rect 384188 566273 384230 566509
rect 383910 566241 384230 566273
rect 389840 566829 390160 566861
rect 389840 566593 389882 566829
rect 390118 566593 390160 566829
rect 389840 566509 390160 566593
rect 389840 566273 389882 566509
rect 390118 566273 390160 566509
rect 389840 566241 390160 566273
rect 395771 566829 396091 566861
rect 395771 566593 395813 566829
rect 396049 566593 396091 566829
rect 395771 566509 396091 566593
rect 395771 566273 395813 566509
rect 396049 566273 396091 566509
rect 395771 566241 396091 566273
rect 411910 566829 412230 566861
rect 411910 566593 411952 566829
rect 412188 566593 412230 566829
rect 411910 566509 412230 566593
rect 411910 566273 411952 566509
rect 412188 566273 412230 566509
rect 411910 566241 412230 566273
rect 417840 566829 418160 566861
rect 417840 566593 417882 566829
rect 418118 566593 418160 566829
rect 417840 566509 418160 566593
rect 417840 566273 417882 566509
rect 418118 566273 418160 566509
rect 417840 566241 418160 566273
rect 423771 566829 424091 566861
rect 423771 566593 423813 566829
rect 424049 566593 424091 566829
rect 423771 566509 424091 566593
rect 423771 566273 423813 566509
rect 424049 566273 424091 566509
rect 423771 566241 424091 566273
rect 439910 566829 440230 566861
rect 439910 566593 439952 566829
rect 440188 566593 440230 566829
rect 439910 566509 440230 566593
rect 439910 566273 439952 566509
rect 440188 566273 440230 566509
rect 439910 566241 440230 566273
rect 445840 566829 446160 566861
rect 445840 566593 445882 566829
rect 446118 566593 446160 566829
rect 445840 566509 446160 566593
rect 445840 566273 445882 566509
rect 446118 566273 446160 566509
rect 445840 566241 446160 566273
rect 451771 566829 452091 566861
rect 451771 566593 451813 566829
rect 452049 566593 452091 566829
rect 451771 566509 452091 566593
rect 451771 566273 451813 566509
rect 452049 566273 452091 566509
rect 451771 566241 452091 566273
rect 467910 566829 468230 566861
rect 467910 566593 467952 566829
rect 468188 566593 468230 566829
rect 467910 566509 468230 566593
rect 467910 566273 467952 566509
rect 468188 566273 468230 566509
rect 467910 566241 468230 566273
rect 473840 566829 474160 566861
rect 473840 566593 473882 566829
rect 474118 566593 474160 566829
rect 473840 566509 474160 566593
rect 473840 566273 473882 566509
rect 474118 566273 474160 566509
rect 473840 566241 474160 566273
rect 479771 566829 480091 566861
rect 479771 566593 479813 566829
rect 480049 566593 480091 566829
rect 479771 566509 480091 566593
rect 479771 566273 479813 566509
rect 480049 566273 480091 566509
rect 479771 566241 480091 566273
rect 495910 566829 496230 566861
rect 495910 566593 495952 566829
rect 496188 566593 496230 566829
rect 495910 566509 496230 566593
rect 495910 566273 495952 566509
rect 496188 566273 496230 566509
rect 495910 566241 496230 566273
rect 501840 566829 502160 566861
rect 501840 566593 501882 566829
rect 502118 566593 502160 566829
rect 501840 566509 502160 566593
rect 501840 566273 501882 566509
rect 502118 566273 502160 566509
rect 501840 566241 502160 566273
rect 507771 566829 508091 566861
rect 507771 566593 507813 566829
rect 508049 566593 508091 566829
rect 507771 566509 508091 566593
rect 507771 566273 507813 566509
rect 508049 566273 508091 566509
rect 507771 566241 508091 566273
rect 523910 566829 524230 566861
rect 523910 566593 523952 566829
rect 524188 566593 524230 566829
rect 523910 566509 524230 566593
rect 523910 566273 523952 566509
rect 524188 566273 524230 566509
rect 523910 566241 524230 566273
rect 529840 566829 530160 566861
rect 529840 566593 529882 566829
rect 530118 566593 530160 566829
rect 529840 566509 530160 566593
rect 529840 566273 529882 566509
rect 530118 566273 530160 566509
rect 529840 566241 530160 566273
rect 535771 566829 536091 566861
rect 535771 566593 535813 566829
rect 536049 566593 536091 566829
rect 535771 566509 536091 566593
rect 535771 566273 535813 566509
rect 536049 566273 536091 566509
rect 535771 566241 536091 566273
rect 551910 566829 552230 566861
rect 551910 566593 551952 566829
rect 552188 566593 552230 566829
rect 551910 566509 552230 566593
rect 551910 566273 551952 566509
rect 552188 566273 552230 566509
rect 551910 566241 552230 566273
rect 557840 566829 558160 566861
rect 557840 566593 557882 566829
rect 558118 566593 558160 566829
rect 557840 566509 558160 566593
rect 557840 566273 557882 566509
rect 558118 566273 558160 566509
rect 557840 566241 558160 566273
rect 563771 566829 564091 566861
rect 563771 566593 563813 566829
rect 564049 566593 564091 566829
rect 563771 566509 564091 566593
rect 563771 566273 563813 566509
rect 564049 566273 564091 566509
rect 563771 566241 564091 566273
rect 573494 566829 574114 593273
rect 573494 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 574114 566829
rect 573494 566509 574114 566593
rect 573494 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 574114 566509
rect 22874 563454 23194 563486
rect 22874 563218 22916 563454
rect 23152 563218 23194 563454
rect 22874 563134 23194 563218
rect 22874 562898 22916 563134
rect 23152 562898 23194 563134
rect 22874 562866 23194 562898
rect 28805 563454 29125 563486
rect 28805 563218 28847 563454
rect 29083 563218 29125 563454
rect 28805 563134 29125 563218
rect 28805 562898 28847 563134
rect 29083 562898 29125 563134
rect 28805 562866 29125 562898
rect 50874 563454 51194 563486
rect 50874 563218 50916 563454
rect 51152 563218 51194 563454
rect 50874 563134 51194 563218
rect 50874 562898 50916 563134
rect 51152 562898 51194 563134
rect 50874 562866 51194 562898
rect 56805 563454 57125 563486
rect 56805 563218 56847 563454
rect 57083 563218 57125 563454
rect 56805 563134 57125 563218
rect 56805 562898 56847 563134
rect 57083 562898 57125 563134
rect 56805 562866 57125 562898
rect 78874 563454 79194 563486
rect 78874 563218 78916 563454
rect 79152 563218 79194 563454
rect 78874 563134 79194 563218
rect 78874 562898 78916 563134
rect 79152 562898 79194 563134
rect 78874 562866 79194 562898
rect 84805 563454 85125 563486
rect 84805 563218 84847 563454
rect 85083 563218 85125 563454
rect 84805 563134 85125 563218
rect 84805 562898 84847 563134
rect 85083 562898 85125 563134
rect 84805 562866 85125 562898
rect 106874 563454 107194 563486
rect 106874 563218 106916 563454
rect 107152 563218 107194 563454
rect 106874 563134 107194 563218
rect 106874 562898 106916 563134
rect 107152 562898 107194 563134
rect 106874 562866 107194 562898
rect 112805 563454 113125 563486
rect 112805 563218 112847 563454
rect 113083 563218 113125 563454
rect 112805 563134 113125 563218
rect 112805 562898 112847 563134
rect 113083 562898 113125 563134
rect 112805 562866 113125 562898
rect 134874 563454 135194 563486
rect 134874 563218 134916 563454
rect 135152 563218 135194 563454
rect 134874 563134 135194 563218
rect 134874 562898 134916 563134
rect 135152 562898 135194 563134
rect 134874 562866 135194 562898
rect 140805 563454 141125 563486
rect 140805 563218 140847 563454
rect 141083 563218 141125 563454
rect 140805 563134 141125 563218
rect 140805 562898 140847 563134
rect 141083 562898 141125 563134
rect 140805 562866 141125 562898
rect 162874 563454 163194 563486
rect 162874 563218 162916 563454
rect 163152 563218 163194 563454
rect 162874 563134 163194 563218
rect 162874 562898 162916 563134
rect 163152 562898 163194 563134
rect 162874 562866 163194 562898
rect 168805 563454 169125 563486
rect 168805 563218 168847 563454
rect 169083 563218 169125 563454
rect 168805 563134 169125 563218
rect 168805 562898 168847 563134
rect 169083 562898 169125 563134
rect 168805 562866 169125 562898
rect 190874 563454 191194 563486
rect 190874 563218 190916 563454
rect 191152 563218 191194 563454
rect 190874 563134 191194 563218
rect 190874 562898 190916 563134
rect 191152 562898 191194 563134
rect 190874 562866 191194 562898
rect 196805 563454 197125 563486
rect 196805 563218 196847 563454
rect 197083 563218 197125 563454
rect 196805 563134 197125 563218
rect 196805 562898 196847 563134
rect 197083 562898 197125 563134
rect 196805 562866 197125 562898
rect 218874 563454 219194 563486
rect 218874 563218 218916 563454
rect 219152 563218 219194 563454
rect 218874 563134 219194 563218
rect 218874 562898 218916 563134
rect 219152 562898 219194 563134
rect 218874 562866 219194 562898
rect 224805 563454 225125 563486
rect 224805 563218 224847 563454
rect 225083 563218 225125 563454
rect 224805 563134 225125 563218
rect 224805 562898 224847 563134
rect 225083 562898 225125 563134
rect 224805 562866 225125 562898
rect 246874 563454 247194 563486
rect 246874 563218 246916 563454
rect 247152 563218 247194 563454
rect 246874 563134 247194 563218
rect 246874 562898 246916 563134
rect 247152 562898 247194 563134
rect 246874 562866 247194 562898
rect 252805 563454 253125 563486
rect 252805 563218 252847 563454
rect 253083 563218 253125 563454
rect 252805 563134 253125 563218
rect 252805 562898 252847 563134
rect 253083 562898 253125 563134
rect 252805 562866 253125 562898
rect 274874 563454 275194 563486
rect 274874 563218 274916 563454
rect 275152 563218 275194 563454
rect 274874 563134 275194 563218
rect 274874 562898 274916 563134
rect 275152 562898 275194 563134
rect 274874 562866 275194 562898
rect 280805 563454 281125 563486
rect 280805 563218 280847 563454
rect 281083 563218 281125 563454
rect 280805 563134 281125 563218
rect 280805 562898 280847 563134
rect 281083 562898 281125 563134
rect 280805 562866 281125 562898
rect 302874 563454 303194 563486
rect 302874 563218 302916 563454
rect 303152 563218 303194 563454
rect 302874 563134 303194 563218
rect 302874 562898 302916 563134
rect 303152 562898 303194 563134
rect 302874 562866 303194 562898
rect 308805 563454 309125 563486
rect 308805 563218 308847 563454
rect 309083 563218 309125 563454
rect 308805 563134 309125 563218
rect 308805 562898 308847 563134
rect 309083 562898 309125 563134
rect 308805 562866 309125 562898
rect 330874 563454 331194 563486
rect 330874 563218 330916 563454
rect 331152 563218 331194 563454
rect 330874 563134 331194 563218
rect 330874 562898 330916 563134
rect 331152 562898 331194 563134
rect 330874 562866 331194 562898
rect 336805 563454 337125 563486
rect 336805 563218 336847 563454
rect 337083 563218 337125 563454
rect 336805 563134 337125 563218
rect 336805 562898 336847 563134
rect 337083 562898 337125 563134
rect 336805 562866 337125 562898
rect 358874 563454 359194 563486
rect 358874 563218 358916 563454
rect 359152 563218 359194 563454
rect 358874 563134 359194 563218
rect 358874 562898 358916 563134
rect 359152 562898 359194 563134
rect 358874 562866 359194 562898
rect 364805 563454 365125 563486
rect 364805 563218 364847 563454
rect 365083 563218 365125 563454
rect 364805 563134 365125 563218
rect 364805 562898 364847 563134
rect 365083 562898 365125 563134
rect 364805 562866 365125 562898
rect 386874 563454 387194 563486
rect 386874 563218 386916 563454
rect 387152 563218 387194 563454
rect 386874 563134 387194 563218
rect 386874 562898 386916 563134
rect 387152 562898 387194 563134
rect 386874 562866 387194 562898
rect 392805 563454 393125 563486
rect 392805 563218 392847 563454
rect 393083 563218 393125 563454
rect 392805 563134 393125 563218
rect 392805 562898 392847 563134
rect 393083 562898 393125 563134
rect 392805 562866 393125 562898
rect 414874 563454 415194 563486
rect 414874 563218 414916 563454
rect 415152 563218 415194 563454
rect 414874 563134 415194 563218
rect 414874 562898 414916 563134
rect 415152 562898 415194 563134
rect 414874 562866 415194 562898
rect 420805 563454 421125 563486
rect 420805 563218 420847 563454
rect 421083 563218 421125 563454
rect 420805 563134 421125 563218
rect 420805 562898 420847 563134
rect 421083 562898 421125 563134
rect 420805 562866 421125 562898
rect 442874 563454 443194 563486
rect 442874 563218 442916 563454
rect 443152 563218 443194 563454
rect 442874 563134 443194 563218
rect 442874 562898 442916 563134
rect 443152 562898 443194 563134
rect 442874 562866 443194 562898
rect 448805 563454 449125 563486
rect 448805 563218 448847 563454
rect 449083 563218 449125 563454
rect 448805 563134 449125 563218
rect 448805 562898 448847 563134
rect 449083 562898 449125 563134
rect 448805 562866 449125 562898
rect 470874 563454 471194 563486
rect 470874 563218 470916 563454
rect 471152 563218 471194 563454
rect 470874 563134 471194 563218
rect 470874 562898 470916 563134
rect 471152 562898 471194 563134
rect 470874 562866 471194 562898
rect 476805 563454 477125 563486
rect 476805 563218 476847 563454
rect 477083 563218 477125 563454
rect 476805 563134 477125 563218
rect 476805 562898 476847 563134
rect 477083 562898 477125 563134
rect 476805 562866 477125 562898
rect 498874 563454 499194 563486
rect 498874 563218 498916 563454
rect 499152 563218 499194 563454
rect 498874 563134 499194 563218
rect 498874 562898 498916 563134
rect 499152 562898 499194 563134
rect 498874 562866 499194 562898
rect 504805 563454 505125 563486
rect 504805 563218 504847 563454
rect 505083 563218 505125 563454
rect 504805 563134 505125 563218
rect 504805 562898 504847 563134
rect 505083 562898 505125 563134
rect 504805 562866 505125 562898
rect 526874 563454 527194 563486
rect 526874 563218 526916 563454
rect 527152 563218 527194 563454
rect 526874 563134 527194 563218
rect 526874 562898 526916 563134
rect 527152 562898 527194 563134
rect 526874 562866 527194 562898
rect 532805 563454 533125 563486
rect 532805 563218 532847 563454
rect 533083 563218 533125 563454
rect 532805 563134 533125 563218
rect 532805 562898 532847 563134
rect 533083 562898 533125 563134
rect 532805 562866 533125 562898
rect 554874 563454 555194 563486
rect 554874 563218 554916 563454
rect 555152 563218 555194 563454
rect 554874 563134 555194 563218
rect 554874 562898 554916 563134
rect 555152 562898 555194 563134
rect 554874 562866 555194 562898
rect 560805 563454 561125 563486
rect 560805 563218 560847 563454
rect 561083 563218 561125 563454
rect 560805 563134 561125 563218
rect 560805 562898 560847 563134
rect 561083 562898 561125 563134
rect 560805 562866 561125 562898
rect -2006 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 -1386 539829
rect -2006 539509 -1386 539593
rect -2006 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 -1386 539509
rect -2006 512829 -1386 539273
rect 19910 539829 20230 539861
rect 19910 539593 19952 539829
rect 20188 539593 20230 539829
rect 19910 539509 20230 539593
rect 19910 539273 19952 539509
rect 20188 539273 20230 539509
rect 19910 539241 20230 539273
rect 25840 539829 26160 539861
rect 25840 539593 25882 539829
rect 26118 539593 26160 539829
rect 25840 539509 26160 539593
rect 25840 539273 25882 539509
rect 26118 539273 26160 539509
rect 25840 539241 26160 539273
rect 31771 539829 32091 539861
rect 31771 539593 31813 539829
rect 32049 539593 32091 539829
rect 31771 539509 32091 539593
rect 31771 539273 31813 539509
rect 32049 539273 32091 539509
rect 31771 539241 32091 539273
rect 47910 539829 48230 539861
rect 47910 539593 47952 539829
rect 48188 539593 48230 539829
rect 47910 539509 48230 539593
rect 47910 539273 47952 539509
rect 48188 539273 48230 539509
rect 47910 539241 48230 539273
rect 53840 539829 54160 539861
rect 53840 539593 53882 539829
rect 54118 539593 54160 539829
rect 53840 539509 54160 539593
rect 53840 539273 53882 539509
rect 54118 539273 54160 539509
rect 53840 539241 54160 539273
rect 59771 539829 60091 539861
rect 59771 539593 59813 539829
rect 60049 539593 60091 539829
rect 59771 539509 60091 539593
rect 59771 539273 59813 539509
rect 60049 539273 60091 539509
rect 59771 539241 60091 539273
rect 75910 539829 76230 539861
rect 75910 539593 75952 539829
rect 76188 539593 76230 539829
rect 75910 539509 76230 539593
rect 75910 539273 75952 539509
rect 76188 539273 76230 539509
rect 75910 539241 76230 539273
rect 81840 539829 82160 539861
rect 81840 539593 81882 539829
rect 82118 539593 82160 539829
rect 81840 539509 82160 539593
rect 81840 539273 81882 539509
rect 82118 539273 82160 539509
rect 81840 539241 82160 539273
rect 87771 539829 88091 539861
rect 87771 539593 87813 539829
rect 88049 539593 88091 539829
rect 87771 539509 88091 539593
rect 87771 539273 87813 539509
rect 88049 539273 88091 539509
rect 87771 539241 88091 539273
rect 103910 539829 104230 539861
rect 103910 539593 103952 539829
rect 104188 539593 104230 539829
rect 103910 539509 104230 539593
rect 103910 539273 103952 539509
rect 104188 539273 104230 539509
rect 103910 539241 104230 539273
rect 109840 539829 110160 539861
rect 109840 539593 109882 539829
rect 110118 539593 110160 539829
rect 109840 539509 110160 539593
rect 109840 539273 109882 539509
rect 110118 539273 110160 539509
rect 109840 539241 110160 539273
rect 115771 539829 116091 539861
rect 115771 539593 115813 539829
rect 116049 539593 116091 539829
rect 115771 539509 116091 539593
rect 115771 539273 115813 539509
rect 116049 539273 116091 539509
rect 115771 539241 116091 539273
rect 131910 539829 132230 539861
rect 131910 539593 131952 539829
rect 132188 539593 132230 539829
rect 131910 539509 132230 539593
rect 131910 539273 131952 539509
rect 132188 539273 132230 539509
rect 131910 539241 132230 539273
rect 137840 539829 138160 539861
rect 137840 539593 137882 539829
rect 138118 539593 138160 539829
rect 137840 539509 138160 539593
rect 137840 539273 137882 539509
rect 138118 539273 138160 539509
rect 137840 539241 138160 539273
rect 143771 539829 144091 539861
rect 143771 539593 143813 539829
rect 144049 539593 144091 539829
rect 143771 539509 144091 539593
rect 143771 539273 143813 539509
rect 144049 539273 144091 539509
rect 143771 539241 144091 539273
rect 159910 539829 160230 539861
rect 159910 539593 159952 539829
rect 160188 539593 160230 539829
rect 159910 539509 160230 539593
rect 159910 539273 159952 539509
rect 160188 539273 160230 539509
rect 159910 539241 160230 539273
rect 165840 539829 166160 539861
rect 165840 539593 165882 539829
rect 166118 539593 166160 539829
rect 165840 539509 166160 539593
rect 165840 539273 165882 539509
rect 166118 539273 166160 539509
rect 165840 539241 166160 539273
rect 171771 539829 172091 539861
rect 171771 539593 171813 539829
rect 172049 539593 172091 539829
rect 171771 539509 172091 539593
rect 171771 539273 171813 539509
rect 172049 539273 172091 539509
rect 171771 539241 172091 539273
rect 187910 539829 188230 539861
rect 187910 539593 187952 539829
rect 188188 539593 188230 539829
rect 187910 539509 188230 539593
rect 187910 539273 187952 539509
rect 188188 539273 188230 539509
rect 187910 539241 188230 539273
rect 193840 539829 194160 539861
rect 193840 539593 193882 539829
rect 194118 539593 194160 539829
rect 193840 539509 194160 539593
rect 193840 539273 193882 539509
rect 194118 539273 194160 539509
rect 193840 539241 194160 539273
rect 199771 539829 200091 539861
rect 199771 539593 199813 539829
rect 200049 539593 200091 539829
rect 199771 539509 200091 539593
rect 199771 539273 199813 539509
rect 200049 539273 200091 539509
rect 199771 539241 200091 539273
rect 215910 539829 216230 539861
rect 215910 539593 215952 539829
rect 216188 539593 216230 539829
rect 215910 539509 216230 539593
rect 215910 539273 215952 539509
rect 216188 539273 216230 539509
rect 215910 539241 216230 539273
rect 221840 539829 222160 539861
rect 221840 539593 221882 539829
rect 222118 539593 222160 539829
rect 221840 539509 222160 539593
rect 221840 539273 221882 539509
rect 222118 539273 222160 539509
rect 221840 539241 222160 539273
rect 227771 539829 228091 539861
rect 227771 539593 227813 539829
rect 228049 539593 228091 539829
rect 227771 539509 228091 539593
rect 227771 539273 227813 539509
rect 228049 539273 228091 539509
rect 227771 539241 228091 539273
rect 243910 539829 244230 539861
rect 243910 539593 243952 539829
rect 244188 539593 244230 539829
rect 243910 539509 244230 539593
rect 243910 539273 243952 539509
rect 244188 539273 244230 539509
rect 243910 539241 244230 539273
rect 249840 539829 250160 539861
rect 249840 539593 249882 539829
rect 250118 539593 250160 539829
rect 249840 539509 250160 539593
rect 249840 539273 249882 539509
rect 250118 539273 250160 539509
rect 249840 539241 250160 539273
rect 255771 539829 256091 539861
rect 255771 539593 255813 539829
rect 256049 539593 256091 539829
rect 255771 539509 256091 539593
rect 255771 539273 255813 539509
rect 256049 539273 256091 539509
rect 255771 539241 256091 539273
rect 271910 539829 272230 539861
rect 271910 539593 271952 539829
rect 272188 539593 272230 539829
rect 271910 539509 272230 539593
rect 271910 539273 271952 539509
rect 272188 539273 272230 539509
rect 271910 539241 272230 539273
rect 277840 539829 278160 539861
rect 277840 539593 277882 539829
rect 278118 539593 278160 539829
rect 277840 539509 278160 539593
rect 277840 539273 277882 539509
rect 278118 539273 278160 539509
rect 277840 539241 278160 539273
rect 283771 539829 284091 539861
rect 283771 539593 283813 539829
rect 284049 539593 284091 539829
rect 283771 539509 284091 539593
rect 283771 539273 283813 539509
rect 284049 539273 284091 539509
rect 283771 539241 284091 539273
rect 299910 539829 300230 539861
rect 299910 539593 299952 539829
rect 300188 539593 300230 539829
rect 299910 539509 300230 539593
rect 299910 539273 299952 539509
rect 300188 539273 300230 539509
rect 299910 539241 300230 539273
rect 305840 539829 306160 539861
rect 305840 539593 305882 539829
rect 306118 539593 306160 539829
rect 305840 539509 306160 539593
rect 305840 539273 305882 539509
rect 306118 539273 306160 539509
rect 305840 539241 306160 539273
rect 311771 539829 312091 539861
rect 311771 539593 311813 539829
rect 312049 539593 312091 539829
rect 311771 539509 312091 539593
rect 311771 539273 311813 539509
rect 312049 539273 312091 539509
rect 311771 539241 312091 539273
rect 327910 539829 328230 539861
rect 327910 539593 327952 539829
rect 328188 539593 328230 539829
rect 327910 539509 328230 539593
rect 327910 539273 327952 539509
rect 328188 539273 328230 539509
rect 327910 539241 328230 539273
rect 333840 539829 334160 539861
rect 333840 539593 333882 539829
rect 334118 539593 334160 539829
rect 333840 539509 334160 539593
rect 333840 539273 333882 539509
rect 334118 539273 334160 539509
rect 333840 539241 334160 539273
rect 339771 539829 340091 539861
rect 339771 539593 339813 539829
rect 340049 539593 340091 539829
rect 339771 539509 340091 539593
rect 339771 539273 339813 539509
rect 340049 539273 340091 539509
rect 339771 539241 340091 539273
rect 355910 539829 356230 539861
rect 355910 539593 355952 539829
rect 356188 539593 356230 539829
rect 355910 539509 356230 539593
rect 355910 539273 355952 539509
rect 356188 539273 356230 539509
rect 355910 539241 356230 539273
rect 361840 539829 362160 539861
rect 361840 539593 361882 539829
rect 362118 539593 362160 539829
rect 361840 539509 362160 539593
rect 361840 539273 361882 539509
rect 362118 539273 362160 539509
rect 361840 539241 362160 539273
rect 367771 539829 368091 539861
rect 367771 539593 367813 539829
rect 368049 539593 368091 539829
rect 367771 539509 368091 539593
rect 367771 539273 367813 539509
rect 368049 539273 368091 539509
rect 367771 539241 368091 539273
rect 383910 539829 384230 539861
rect 383910 539593 383952 539829
rect 384188 539593 384230 539829
rect 383910 539509 384230 539593
rect 383910 539273 383952 539509
rect 384188 539273 384230 539509
rect 383910 539241 384230 539273
rect 389840 539829 390160 539861
rect 389840 539593 389882 539829
rect 390118 539593 390160 539829
rect 389840 539509 390160 539593
rect 389840 539273 389882 539509
rect 390118 539273 390160 539509
rect 389840 539241 390160 539273
rect 395771 539829 396091 539861
rect 395771 539593 395813 539829
rect 396049 539593 396091 539829
rect 395771 539509 396091 539593
rect 395771 539273 395813 539509
rect 396049 539273 396091 539509
rect 395771 539241 396091 539273
rect 411910 539829 412230 539861
rect 411910 539593 411952 539829
rect 412188 539593 412230 539829
rect 411910 539509 412230 539593
rect 411910 539273 411952 539509
rect 412188 539273 412230 539509
rect 411910 539241 412230 539273
rect 417840 539829 418160 539861
rect 417840 539593 417882 539829
rect 418118 539593 418160 539829
rect 417840 539509 418160 539593
rect 417840 539273 417882 539509
rect 418118 539273 418160 539509
rect 417840 539241 418160 539273
rect 423771 539829 424091 539861
rect 423771 539593 423813 539829
rect 424049 539593 424091 539829
rect 423771 539509 424091 539593
rect 423771 539273 423813 539509
rect 424049 539273 424091 539509
rect 423771 539241 424091 539273
rect 439910 539829 440230 539861
rect 439910 539593 439952 539829
rect 440188 539593 440230 539829
rect 439910 539509 440230 539593
rect 439910 539273 439952 539509
rect 440188 539273 440230 539509
rect 439910 539241 440230 539273
rect 445840 539829 446160 539861
rect 445840 539593 445882 539829
rect 446118 539593 446160 539829
rect 445840 539509 446160 539593
rect 445840 539273 445882 539509
rect 446118 539273 446160 539509
rect 445840 539241 446160 539273
rect 451771 539829 452091 539861
rect 451771 539593 451813 539829
rect 452049 539593 452091 539829
rect 451771 539509 452091 539593
rect 451771 539273 451813 539509
rect 452049 539273 452091 539509
rect 451771 539241 452091 539273
rect 467910 539829 468230 539861
rect 467910 539593 467952 539829
rect 468188 539593 468230 539829
rect 467910 539509 468230 539593
rect 467910 539273 467952 539509
rect 468188 539273 468230 539509
rect 467910 539241 468230 539273
rect 473840 539829 474160 539861
rect 473840 539593 473882 539829
rect 474118 539593 474160 539829
rect 473840 539509 474160 539593
rect 473840 539273 473882 539509
rect 474118 539273 474160 539509
rect 473840 539241 474160 539273
rect 479771 539829 480091 539861
rect 479771 539593 479813 539829
rect 480049 539593 480091 539829
rect 479771 539509 480091 539593
rect 479771 539273 479813 539509
rect 480049 539273 480091 539509
rect 479771 539241 480091 539273
rect 495910 539829 496230 539861
rect 495910 539593 495952 539829
rect 496188 539593 496230 539829
rect 495910 539509 496230 539593
rect 495910 539273 495952 539509
rect 496188 539273 496230 539509
rect 495910 539241 496230 539273
rect 501840 539829 502160 539861
rect 501840 539593 501882 539829
rect 502118 539593 502160 539829
rect 501840 539509 502160 539593
rect 501840 539273 501882 539509
rect 502118 539273 502160 539509
rect 501840 539241 502160 539273
rect 507771 539829 508091 539861
rect 507771 539593 507813 539829
rect 508049 539593 508091 539829
rect 507771 539509 508091 539593
rect 507771 539273 507813 539509
rect 508049 539273 508091 539509
rect 507771 539241 508091 539273
rect 523910 539829 524230 539861
rect 523910 539593 523952 539829
rect 524188 539593 524230 539829
rect 523910 539509 524230 539593
rect 523910 539273 523952 539509
rect 524188 539273 524230 539509
rect 523910 539241 524230 539273
rect 529840 539829 530160 539861
rect 529840 539593 529882 539829
rect 530118 539593 530160 539829
rect 529840 539509 530160 539593
rect 529840 539273 529882 539509
rect 530118 539273 530160 539509
rect 529840 539241 530160 539273
rect 535771 539829 536091 539861
rect 535771 539593 535813 539829
rect 536049 539593 536091 539829
rect 535771 539509 536091 539593
rect 535771 539273 535813 539509
rect 536049 539273 536091 539509
rect 535771 539241 536091 539273
rect 551910 539829 552230 539861
rect 551910 539593 551952 539829
rect 552188 539593 552230 539829
rect 551910 539509 552230 539593
rect 551910 539273 551952 539509
rect 552188 539273 552230 539509
rect 551910 539241 552230 539273
rect 557840 539829 558160 539861
rect 557840 539593 557882 539829
rect 558118 539593 558160 539829
rect 557840 539509 558160 539593
rect 557840 539273 557882 539509
rect 558118 539273 558160 539509
rect 557840 539241 558160 539273
rect 563771 539829 564091 539861
rect 563771 539593 563813 539829
rect 564049 539593 564091 539829
rect 563771 539509 564091 539593
rect 563771 539273 563813 539509
rect 564049 539273 564091 539509
rect 563771 539241 564091 539273
rect 573494 539829 574114 566273
rect 573494 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 574114 539829
rect 573494 539509 574114 539593
rect 573494 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 574114 539509
rect 22874 536454 23194 536486
rect 22874 536218 22916 536454
rect 23152 536218 23194 536454
rect 22874 536134 23194 536218
rect 22874 535898 22916 536134
rect 23152 535898 23194 536134
rect 22874 535866 23194 535898
rect 28805 536454 29125 536486
rect 28805 536218 28847 536454
rect 29083 536218 29125 536454
rect 28805 536134 29125 536218
rect 28805 535898 28847 536134
rect 29083 535898 29125 536134
rect 28805 535866 29125 535898
rect 50874 536454 51194 536486
rect 50874 536218 50916 536454
rect 51152 536218 51194 536454
rect 50874 536134 51194 536218
rect 50874 535898 50916 536134
rect 51152 535898 51194 536134
rect 50874 535866 51194 535898
rect 56805 536454 57125 536486
rect 56805 536218 56847 536454
rect 57083 536218 57125 536454
rect 56805 536134 57125 536218
rect 56805 535898 56847 536134
rect 57083 535898 57125 536134
rect 56805 535866 57125 535898
rect 78874 536454 79194 536486
rect 78874 536218 78916 536454
rect 79152 536218 79194 536454
rect 78874 536134 79194 536218
rect 78874 535898 78916 536134
rect 79152 535898 79194 536134
rect 78874 535866 79194 535898
rect 84805 536454 85125 536486
rect 84805 536218 84847 536454
rect 85083 536218 85125 536454
rect 84805 536134 85125 536218
rect 84805 535898 84847 536134
rect 85083 535898 85125 536134
rect 84805 535866 85125 535898
rect 106874 536454 107194 536486
rect 106874 536218 106916 536454
rect 107152 536218 107194 536454
rect 106874 536134 107194 536218
rect 106874 535898 106916 536134
rect 107152 535898 107194 536134
rect 106874 535866 107194 535898
rect 112805 536454 113125 536486
rect 112805 536218 112847 536454
rect 113083 536218 113125 536454
rect 112805 536134 113125 536218
rect 112805 535898 112847 536134
rect 113083 535898 113125 536134
rect 112805 535866 113125 535898
rect 134874 536454 135194 536486
rect 134874 536218 134916 536454
rect 135152 536218 135194 536454
rect 134874 536134 135194 536218
rect 134874 535898 134916 536134
rect 135152 535898 135194 536134
rect 134874 535866 135194 535898
rect 140805 536454 141125 536486
rect 140805 536218 140847 536454
rect 141083 536218 141125 536454
rect 140805 536134 141125 536218
rect 140805 535898 140847 536134
rect 141083 535898 141125 536134
rect 140805 535866 141125 535898
rect 162874 536454 163194 536486
rect 162874 536218 162916 536454
rect 163152 536218 163194 536454
rect 162874 536134 163194 536218
rect 162874 535898 162916 536134
rect 163152 535898 163194 536134
rect 162874 535866 163194 535898
rect 168805 536454 169125 536486
rect 168805 536218 168847 536454
rect 169083 536218 169125 536454
rect 168805 536134 169125 536218
rect 168805 535898 168847 536134
rect 169083 535898 169125 536134
rect 168805 535866 169125 535898
rect 190874 536454 191194 536486
rect 190874 536218 190916 536454
rect 191152 536218 191194 536454
rect 190874 536134 191194 536218
rect 190874 535898 190916 536134
rect 191152 535898 191194 536134
rect 190874 535866 191194 535898
rect 196805 536454 197125 536486
rect 196805 536218 196847 536454
rect 197083 536218 197125 536454
rect 196805 536134 197125 536218
rect 196805 535898 196847 536134
rect 197083 535898 197125 536134
rect 196805 535866 197125 535898
rect 218874 536454 219194 536486
rect 218874 536218 218916 536454
rect 219152 536218 219194 536454
rect 218874 536134 219194 536218
rect 218874 535898 218916 536134
rect 219152 535898 219194 536134
rect 218874 535866 219194 535898
rect 224805 536454 225125 536486
rect 224805 536218 224847 536454
rect 225083 536218 225125 536454
rect 224805 536134 225125 536218
rect 224805 535898 224847 536134
rect 225083 535898 225125 536134
rect 224805 535866 225125 535898
rect 246874 536454 247194 536486
rect 246874 536218 246916 536454
rect 247152 536218 247194 536454
rect 246874 536134 247194 536218
rect 246874 535898 246916 536134
rect 247152 535898 247194 536134
rect 246874 535866 247194 535898
rect 252805 536454 253125 536486
rect 252805 536218 252847 536454
rect 253083 536218 253125 536454
rect 252805 536134 253125 536218
rect 252805 535898 252847 536134
rect 253083 535898 253125 536134
rect 252805 535866 253125 535898
rect 274874 536454 275194 536486
rect 274874 536218 274916 536454
rect 275152 536218 275194 536454
rect 274874 536134 275194 536218
rect 274874 535898 274916 536134
rect 275152 535898 275194 536134
rect 274874 535866 275194 535898
rect 280805 536454 281125 536486
rect 280805 536218 280847 536454
rect 281083 536218 281125 536454
rect 280805 536134 281125 536218
rect 280805 535898 280847 536134
rect 281083 535898 281125 536134
rect 280805 535866 281125 535898
rect 302874 536454 303194 536486
rect 302874 536218 302916 536454
rect 303152 536218 303194 536454
rect 302874 536134 303194 536218
rect 302874 535898 302916 536134
rect 303152 535898 303194 536134
rect 302874 535866 303194 535898
rect 308805 536454 309125 536486
rect 308805 536218 308847 536454
rect 309083 536218 309125 536454
rect 308805 536134 309125 536218
rect 308805 535898 308847 536134
rect 309083 535898 309125 536134
rect 308805 535866 309125 535898
rect 330874 536454 331194 536486
rect 330874 536218 330916 536454
rect 331152 536218 331194 536454
rect 330874 536134 331194 536218
rect 330874 535898 330916 536134
rect 331152 535898 331194 536134
rect 330874 535866 331194 535898
rect 336805 536454 337125 536486
rect 336805 536218 336847 536454
rect 337083 536218 337125 536454
rect 336805 536134 337125 536218
rect 336805 535898 336847 536134
rect 337083 535898 337125 536134
rect 336805 535866 337125 535898
rect 358874 536454 359194 536486
rect 358874 536218 358916 536454
rect 359152 536218 359194 536454
rect 358874 536134 359194 536218
rect 358874 535898 358916 536134
rect 359152 535898 359194 536134
rect 358874 535866 359194 535898
rect 364805 536454 365125 536486
rect 364805 536218 364847 536454
rect 365083 536218 365125 536454
rect 364805 536134 365125 536218
rect 364805 535898 364847 536134
rect 365083 535898 365125 536134
rect 364805 535866 365125 535898
rect 386874 536454 387194 536486
rect 386874 536218 386916 536454
rect 387152 536218 387194 536454
rect 386874 536134 387194 536218
rect 386874 535898 386916 536134
rect 387152 535898 387194 536134
rect 386874 535866 387194 535898
rect 392805 536454 393125 536486
rect 392805 536218 392847 536454
rect 393083 536218 393125 536454
rect 392805 536134 393125 536218
rect 392805 535898 392847 536134
rect 393083 535898 393125 536134
rect 392805 535866 393125 535898
rect 414874 536454 415194 536486
rect 414874 536218 414916 536454
rect 415152 536218 415194 536454
rect 414874 536134 415194 536218
rect 414874 535898 414916 536134
rect 415152 535898 415194 536134
rect 414874 535866 415194 535898
rect 420805 536454 421125 536486
rect 420805 536218 420847 536454
rect 421083 536218 421125 536454
rect 420805 536134 421125 536218
rect 420805 535898 420847 536134
rect 421083 535898 421125 536134
rect 420805 535866 421125 535898
rect 442874 536454 443194 536486
rect 442874 536218 442916 536454
rect 443152 536218 443194 536454
rect 442874 536134 443194 536218
rect 442874 535898 442916 536134
rect 443152 535898 443194 536134
rect 442874 535866 443194 535898
rect 448805 536454 449125 536486
rect 448805 536218 448847 536454
rect 449083 536218 449125 536454
rect 448805 536134 449125 536218
rect 448805 535898 448847 536134
rect 449083 535898 449125 536134
rect 448805 535866 449125 535898
rect 470874 536454 471194 536486
rect 470874 536218 470916 536454
rect 471152 536218 471194 536454
rect 470874 536134 471194 536218
rect 470874 535898 470916 536134
rect 471152 535898 471194 536134
rect 470874 535866 471194 535898
rect 476805 536454 477125 536486
rect 476805 536218 476847 536454
rect 477083 536218 477125 536454
rect 476805 536134 477125 536218
rect 476805 535898 476847 536134
rect 477083 535898 477125 536134
rect 476805 535866 477125 535898
rect 498874 536454 499194 536486
rect 498874 536218 498916 536454
rect 499152 536218 499194 536454
rect 498874 536134 499194 536218
rect 498874 535898 498916 536134
rect 499152 535898 499194 536134
rect 498874 535866 499194 535898
rect 504805 536454 505125 536486
rect 504805 536218 504847 536454
rect 505083 536218 505125 536454
rect 504805 536134 505125 536218
rect 504805 535898 504847 536134
rect 505083 535898 505125 536134
rect 504805 535866 505125 535898
rect 526874 536454 527194 536486
rect 526874 536218 526916 536454
rect 527152 536218 527194 536454
rect 526874 536134 527194 536218
rect 526874 535898 526916 536134
rect 527152 535898 527194 536134
rect 526874 535866 527194 535898
rect 532805 536454 533125 536486
rect 532805 536218 532847 536454
rect 533083 536218 533125 536454
rect 532805 536134 533125 536218
rect 532805 535898 532847 536134
rect 533083 535898 533125 536134
rect 532805 535866 533125 535898
rect 554874 536454 555194 536486
rect 554874 536218 554916 536454
rect 555152 536218 555194 536454
rect 554874 536134 555194 536218
rect 554874 535898 554916 536134
rect 555152 535898 555194 536134
rect 554874 535866 555194 535898
rect 560805 536454 561125 536486
rect 560805 536218 560847 536454
rect 561083 536218 561125 536454
rect 560805 536134 561125 536218
rect 560805 535898 560847 536134
rect 561083 535898 561125 536134
rect 560805 535866 561125 535898
rect -2006 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 -1386 512829
rect -2006 512509 -1386 512593
rect -2006 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 -1386 512509
rect -2006 485829 -1386 512273
rect 19910 512829 20230 512861
rect 19910 512593 19952 512829
rect 20188 512593 20230 512829
rect 19910 512509 20230 512593
rect 19910 512273 19952 512509
rect 20188 512273 20230 512509
rect 19910 512241 20230 512273
rect 25840 512829 26160 512861
rect 25840 512593 25882 512829
rect 26118 512593 26160 512829
rect 25840 512509 26160 512593
rect 25840 512273 25882 512509
rect 26118 512273 26160 512509
rect 25840 512241 26160 512273
rect 31771 512829 32091 512861
rect 31771 512593 31813 512829
rect 32049 512593 32091 512829
rect 31771 512509 32091 512593
rect 31771 512273 31813 512509
rect 32049 512273 32091 512509
rect 31771 512241 32091 512273
rect 47910 512829 48230 512861
rect 47910 512593 47952 512829
rect 48188 512593 48230 512829
rect 47910 512509 48230 512593
rect 47910 512273 47952 512509
rect 48188 512273 48230 512509
rect 47910 512241 48230 512273
rect 53840 512829 54160 512861
rect 53840 512593 53882 512829
rect 54118 512593 54160 512829
rect 53840 512509 54160 512593
rect 53840 512273 53882 512509
rect 54118 512273 54160 512509
rect 53840 512241 54160 512273
rect 59771 512829 60091 512861
rect 59771 512593 59813 512829
rect 60049 512593 60091 512829
rect 59771 512509 60091 512593
rect 59771 512273 59813 512509
rect 60049 512273 60091 512509
rect 59771 512241 60091 512273
rect 75910 512829 76230 512861
rect 75910 512593 75952 512829
rect 76188 512593 76230 512829
rect 75910 512509 76230 512593
rect 75910 512273 75952 512509
rect 76188 512273 76230 512509
rect 75910 512241 76230 512273
rect 81840 512829 82160 512861
rect 81840 512593 81882 512829
rect 82118 512593 82160 512829
rect 81840 512509 82160 512593
rect 81840 512273 81882 512509
rect 82118 512273 82160 512509
rect 81840 512241 82160 512273
rect 87771 512829 88091 512861
rect 87771 512593 87813 512829
rect 88049 512593 88091 512829
rect 87771 512509 88091 512593
rect 87771 512273 87813 512509
rect 88049 512273 88091 512509
rect 87771 512241 88091 512273
rect 103910 512829 104230 512861
rect 103910 512593 103952 512829
rect 104188 512593 104230 512829
rect 103910 512509 104230 512593
rect 103910 512273 103952 512509
rect 104188 512273 104230 512509
rect 103910 512241 104230 512273
rect 109840 512829 110160 512861
rect 109840 512593 109882 512829
rect 110118 512593 110160 512829
rect 109840 512509 110160 512593
rect 109840 512273 109882 512509
rect 110118 512273 110160 512509
rect 109840 512241 110160 512273
rect 115771 512829 116091 512861
rect 115771 512593 115813 512829
rect 116049 512593 116091 512829
rect 115771 512509 116091 512593
rect 115771 512273 115813 512509
rect 116049 512273 116091 512509
rect 115771 512241 116091 512273
rect 131910 512829 132230 512861
rect 131910 512593 131952 512829
rect 132188 512593 132230 512829
rect 131910 512509 132230 512593
rect 131910 512273 131952 512509
rect 132188 512273 132230 512509
rect 131910 512241 132230 512273
rect 137840 512829 138160 512861
rect 137840 512593 137882 512829
rect 138118 512593 138160 512829
rect 137840 512509 138160 512593
rect 137840 512273 137882 512509
rect 138118 512273 138160 512509
rect 137840 512241 138160 512273
rect 143771 512829 144091 512861
rect 143771 512593 143813 512829
rect 144049 512593 144091 512829
rect 143771 512509 144091 512593
rect 143771 512273 143813 512509
rect 144049 512273 144091 512509
rect 143771 512241 144091 512273
rect 159910 512829 160230 512861
rect 159910 512593 159952 512829
rect 160188 512593 160230 512829
rect 159910 512509 160230 512593
rect 159910 512273 159952 512509
rect 160188 512273 160230 512509
rect 159910 512241 160230 512273
rect 165840 512829 166160 512861
rect 165840 512593 165882 512829
rect 166118 512593 166160 512829
rect 165840 512509 166160 512593
rect 165840 512273 165882 512509
rect 166118 512273 166160 512509
rect 165840 512241 166160 512273
rect 171771 512829 172091 512861
rect 171771 512593 171813 512829
rect 172049 512593 172091 512829
rect 171771 512509 172091 512593
rect 171771 512273 171813 512509
rect 172049 512273 172091 512509
rect 171771 512241 172091 512273
rect 187910 512829 188230 512861
rect 187910 512593 187952 512829
rect 188188 512593 188230 512829
rect 187910 512509 188230 512593
rect 187910 512273 187952 512509
rect 188188 512273 188230 512509
rect 187910 512241 188230 512273
rect 193840 512829 194160 512861
rect 193840 512593 193882 512829
rect 194118 512593 194160 512829
rect 193840 512509 194160 512593
rect 193840 512273 193882 512509
rect 194118 512273 194160 512509
rect 193840 512241 194160 512273
rect 199771 512829 200091 512861
rect 199771 512593 199813 512829
rect 200049 512593 200091 512829
rect 199771 512509 200091 512593
rect 199771 512273 199813 512509
rect 200049 512273 200091 512509
rect 199771 512241 200091 512273
rect 215910 512829 216230 512861
rect 215910 512593 215952 512829
rect 216188 512593 216230 512829
rect 215910 512509 216230 512593
rect 215910 512273 215952 512509
rect 216188 512273 216230 512509
rect 215910 512241 216230 512273
rect 221840 512829 222160 512861
rect 221840 512593 221882 512829
rect 222118 512593 222160 512829
rect 221840 512509 222160 512593
rect 221840 512273 221882 512509
rect 222118 512273 222160 512509
rect 221840 512241 222160 512273
rect 227771 512829 228091 512861
rect 227771 512593 227813 512829
rect 228049 512593 228091 512829
rect 227771 512509 228091 512593
rect 227771 512273 227813 512509
rect 228049 512273 228091 512509
rect 227771 512241 228091 512273
rect 243910 512829 244230 512861
rect 243910 512593 243952 512829
rect 244188 512593 244230 512829
rect 243910 512509 244230 512593
rect 243910 512273 243952 512509
rect 244188 512273 244230 512509
rect 243910 512241 244230 512273
rect 249840 512829 250160 512861
rect 249840 512593 249882 512829
rect 250118 512593 250160 512829
rect 249840 512509 250160 512593
rect 249840 512273 249882 512509
rect 250118 512273 250160 512509
rect 249840 512241 250160 512273
rect 255771 512829 256091 512861
rect 255771 512593 255813 512829
rect 256049 512593 256091 512829
rect 255771 512509 256091 512593
rect 255771 512273 255813 512509
rect 256049 512273 256091 512509
rect 255771 512241 256091 512273
rect 271910 512829 272230 512861
rect 271910 512593 271952 512829
rect 272188 512593 272230 512829
rect 271910 512509 272230 512593
rect 271910 512273 271952 512509
rect 272188 512273 272230 512509
rect 271910 512241 272230 512273
rect 277840 512829 278160 512861
rect 277840 512593 277882 512829
rect 278118 512593 278160 512829
rect 277840 512509 278160 512593
rect 277840 512273 277882 512509
rect 278118 512273 278160 512509
rect 277840 512241 278160 512273
rect 283771 512829 284091 512861
rect 283771 512593 283813 512829
rect 284049 512593 284091 512829
rect 283771 512509 284091 512593
rect 283771 512273 283813 512509
rect 284049 512273 284091 512509
rect 283771 512241 284091 512273
rect 299910 512829 300230 512861
rect 299910 512593 299952 512829
rect 300188 512593 300230 512829
rect 299910 512509 300230 512593
rect 299910 512273 299952 512509
rect 300188 512273 300230 512509
rect 299910 512241 300230 512273
rect 305840 512829 306160 512861
rect 305840 512593 305882 512829
rect 306118 512593 306160 512829
rect 305840 512509 306160 512593
rect 305840 512273 305882 512509
rect 306118 512273 306160 512509
rect 305840 512241 306160 512273
rect 311771 512829 312091 512861
rect 311771 512593 311813 512829
rect 312049 512593 312091 512829
rect 311771 512509 312091 512593
rect 311771 512273 311813 512509
rect 312049 512273 312091 512509
rect 311771 512241 312091 512273
rect 327910 512829 328230 512861
rect 327910 512593 327952 512829
rect 328188 512593 328230 512829
rect 327910 512509 328230 512593
rect 327910 512273 327952 512509
rect 328188 512273 328230 512509
rect 327910 512241 328230 512273
rect 333840 512829 334160 512861
rect 333840 512593 333882 512829
rect 334118 512593 334160 512829
rect 333840 512509 334160 512593
rect 333840 512273 333882 512509
rect 334118 512273 334160 512509
rect 333840 512241 334160 512273
rect 339771 512829 340091 512861
rect 339771 512593 339813 512829
rect 340049 512593 340091 512829
rect 339771 512509 340091 512593
rect 339771 512273 339813 512509
rect 340049 512273 340091 512509
rect 339771 512241 340091 512273
rect 355910 512829 356230 512861
rect 355910 512593 355952 512829
rect 356188 512593 356230 512829
rect 355910 512509 356230 512593
rect 355910 512273 355952 512509
rect 356188 512273 356230 512509
rect 355910 512241 356230 512273
rect 361840 512829 362160 512861
rect 361840 512593 361882 512829
rect 362118 512593 362160 512829
rect 361840 512509 362160 512593
rect 361840 512273 361882 512509
rect 362118 512273 362160 512509
rect 361840 512241 362160 512273
rect 367771 512829 368091 512861
rect 367771 512593 367813 512829
rect 368049 512593 368091 512829
rect 367771 512509 368091 512593
rect 367771 512273 367813 512509
rect 368049 512273 368091 512509
rect 367771 512241 368091 512273
rect 383910 512829 384230 512861
rect 383910 512593 383952 512829
rect 384188 512593 384230 512829
rect 383910 512509 384230 512593
rect 383910 512273 383952 512509
rect 384188 512273 384230 512509
rect 383910 512241 384230 512273
rect 389840 512829 390160 512861
rect 389840 512593 389882 512829
rect 390118 512593 390160 512829
rect 389840 512509 390160 512593
rect 389840 512273 389882 512509
rect 390118 512273 390160 512509
rect 389840 512241 390160 512273
rect 395771 512829 396091 512861
rect 395771 512593 395813 512829
rect 396049 512593 396091 512829
rect 395771 512509 396091 512593
rect 395771 512273 395813 512509
rect 396049 512273 396091 512509
rect 395771 512241 396091 512273
rect 411910 512829 412230 512861
rect 411910 512593 411952 512829
rect 412188 512593 412230 512829
rect 411910 512509 412230 512593
rect 411910 512273 411952 512509
rect 412188 512273 412230 512509
rect 411910 512241 412230 512273
rect 417840 512829 418160 512861
rect 417840 512593 417882 512829
rect 418118 512593 418160 512829
rect 417840 512509 418160 512593
rect 417840 512273 417882 512509
rect 418118 512273 418160 512509
rect 417840 512241 418160 512273
rect 423771 512829 424091 512861
rect 423771 512593 423813 512829
rect 424049 512593 424091 512829
rect 423771 512509 424091 512593
rect 423771 512273 423813 512509
rect 424049 512273 424091 512509
rect 423771 512241 424091 512273
rect 439910 512829 440230 512861
rect 439910 512593 439952 512829
rect 440188 512593 440230 512829
rect 439910 512509 440230 512593
rect 439910 512273 439952 512509
rect 440188 512273 440230 512509
rect 439910 512241 440230 512273
rect 445840 512829 446160 512861
rect 445840 512593 445882 512829
rect 446118 512593 446160 512829
rect 445840 512509 446160 512593
rect 445840 512273 445882 512509
rect 446118 512273 446160 512509
rect 445840 512241 446160 512273
rect 451771 512829 452091 512861
rect 451771 512593 451813 512829
rect 452049 512593 452091 512829
rect 451771 512509 452091 512593
rect 451771 512273 451813 512509
rect 452049 512273 452091 512509
rect 451771 512241 452091 512273
rect 467910 512829 468230 512861
rect 467910 512593 467952 512829
rect 468188 512593 468230 512829
rect 467910 512509 468230 512593
rect 467910 512273 467952 512509
rect 468188 512273 468230 512509
rect 467910 512241 468230 512273
rect 473840 512829 474160 512861
rect 473840 512593 473882 512829
rect 474118 512593 474160 512829
rect 473840 512509 474160 512593
rect 473840 512273 473882 512509
rect 474118 512273 474160 512509
rect 473840 512241 474160 512273
rect 479771 512829 480091 512861
rect 479771 512593 479813 512829
rect 480049 512593 480091 512829
rect 479771 512509 480091 512593
rect 479771 512273 479813 512509
rect 480049 512273 480091 512509
rect 479771 512241 480091 512273
rect 495910 512829 496230 512861
rect 495910 512593 495952 512829
rect 496188 512593 496230 512829
rect 495910 512509 496230 512593
rect 495910 512273 495952 512509
rect 496188 512273 496230 512509
rect 495910 512241 496230 512273
rect 501840 512829 502160 512861
rect 501840 512593 501882 512829
rect 502118 512593 502160 512829
rect 501840 512509 502160 512593
rect 501840 512273 501882 512509
rect 502118 512273 502160 512509
rect 501840 512241 502160 512273
rect 507771 512829 508091 512861
rect 507771 512593 507813 512829
rect 508049 512593 508091 512829
rect 507771 512509 508091 512593
rect 507771 512273 507813 512509
rect 508049 512273 508091 512509
rect 507771 512241 508091 512273
rect 523910 512829 524230 512861
rect 523910 512593 523952 512829
rect 524188 512593 524230 512829
rect 523910 512509 524230 512593
rect 523910 512273 523952 512509
rect 524188 512273 524230 512509
rect 523910 512241 524230 512273
rect 529840 512829 530160 512861
rect 529840 512593 529882 512829
rect 530118 512593 530160 512829
rect 529840 512509 530160 512593
rect 529840 512273 529882 512509
rect 530118 512273 530160 512509
rect 529840 512241 530160 512273
rect 535771 512829 536091 512861
rect 535771 512593 535813 512829
rect 536049 512593 536091 512829
rect 535771 512509 536091 512593
rect 535771 512273 535813 512509
rect 536049 512273 536091 512509
rect 535771 512241 536091 512273
rect 551910 512829 552230 512861
rect 551910 512593 551952 512829
rect 552188 512593 552230 512829
rect 551910 512509 552230 512593
rect 551910 512273 551952 512509
rect 552188 512273 552230 512509
rect 551910 512241 552230 512273
rect 557840 512829 558160 512861
rect 557840 512593 557882 512829
rect 558118 512593 558160 512829
rect 557840 512509 558160 512593
rect 557840 512273 557882 512509
rect 558118 512273 558160 512509
rect 557840 512241 558160 512273
rect 563771 512829 564091 512861
rect 563771 512593 563813 512829
rect 564049 512593 564091 512829
rect 563771 512509 564091 512593
rect 563771 512273 563813 512509
rect 564049 512273 564091 512509
rect 563771 512241 564091 512273
rect 573494 512829 574114 539273
rect 573494 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 574114 512829
rect 573494 512509 574114 512593
rect 573494 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 574114 512509
rect 22874 509454 23194 509486
rect 22874 509218 22916 509454
rect 23152 509218 23194 509454
rect 22874 509134 23194 509218
rect 22874 508898 22916 509134
rect 23152 508898 23194 509134
rect 22874 508866 23194 508898
rect 28805 509454 29125 509486
rect 28805 509218 28847 509454
rect 29083 509218 29125 509454
rect 28805 509134 29125 509218
rect 28805 508898 28847 509134
rect 29083 508898 29125 509134
rect 28805 508866 29125 508898
rect 50874 509454 51194 509486
rect 50874 509218 50916 509454
rect 51152 509218 51194 509454
rect 50874 509134 51194 509218
rect 50874 508898 50916 509134
rect 51152 508898 51194 509134
rect 50874 508866 51194 508898
rect 56805 509454 57125 509486
rect 56805 509218 56847 509454
rect 57083 509218 57125 509454
rect 56805 509134 57125 509218
rect 56805 508898 56847 509134
rect 57083 508898 57125 509134
rect 56805 508866 57125 508898
rect 78874 509454 79194 509486
rect 78874 509218 78916 509454
rect 79152 509218 79194 509454
rect 78874 509134 79194 509218
rect 78874 508898 78916 509134
rect 79152 508898 79194 509134
rect 78874 508866 79194 508898
rect 84805 509454 85125 509486
rect 84805 509218 84847 509454
rect 85083 509218 85125 509454
rect 84805 509134 85125 509218
rect 84805 508898 84847 509134
rect 85083 508898 85125 509134
rect 84805 508866 85125 508898
rect 106874 509454 107194 509486
rect 106874 509218 106916 509454
rect 107152 509218 107194 509454
rect 106874 509134 107194 509218
rect 106874 508898 106916 509134
rect 107152 508898 107194 509134
rect 106874 508866 107194 508898
rect 112805 509454 113125 509486
rect 112805 509218 112847 509454
rect 113083 509218 113125 509454
rect 112805 509134 113125 509218
rect 112805 508898 112847 509134
rect 113083 508898 113125 509134
rect 112805 508866 113125 508898
rect 134874 509454 135194 509486
rect 134874 509218 134916 509454
rect 135152 509218 135194 509454
rect 134874 509134 135194 509218
rect 134874 508898 134916 509134
rect 135152 508898 135194 509134
rect 134874 508866 135194 508898
rect 140805 509454 141125 509486
rect 140805 509218 140847 509454
rect 141083 509218 141125 509454
rect 140805 509134 141125 509218
rect 140805 508898 140847 509134
rect 141083 508898 141125 509134
rect 140805 508866 141125 508898
rect 162874 509454 163194 509486
rect 162874 509218 162916 509454
rect 163152 509218 163194 509454
rect 162874 509134 163194 509218
rect 162874 508898 162916 509134
rect 163152 508898 163194 509134
rect 162874 508866 163194 508898
rect 168805 509454 169125 509486
rect 168805 509218 168847 509454
rect 169083 509218 169125 509454
rect 168805 509134 169125 509218
rect 168805 508898 168847 509134
rect 169083 508898 169125 509134
rect 168805 508866 169125 508898
rect 190874 509454 191194 509486
rect 190874 509218 190916 509454
rect 191152 509218 191194 509454
rect 190874 509134 191194 509218
rect 190874 508898 190916 509134
rect 191152 508898 191194 509134
rect 190874 508866 191194 508898
rect 196805 509454 197125 509486
rect 196805 509218 196847 509454
rect 197083 509218 197125 509454
rect 196805 509134 197125 509218
rect 196805 508898 196847 509134
rect 197083 508898 197125 509134
rect 196805 508866 197125 508898
rect 218874 509454 219194 509486
rect 218874 509218 218916 509454
rect 219152 509218 219194 509454
rect 218874 509134 219194 509218
rect 218874 508898 218916 509134
rect 219152 508898 219194 509134
rect 218874 508866 219194 508898
rect 224805 509454 225125 509486
rect 224805 509218 224847 509454
rect 225083 509218 225125 509454
rect 224805 509134 225125 509218
rect 224805 508898 224847 509134
rect 225083 508898 225125 509134
rect 224805 508866 225125 508898
rect 246874 509454 247194 509486
rect 246874 509218 246916 509454
rect 247152 509218 247194 509454
rect 246874 509134 247194 509218
rect 246874 508898 246916 509134
rect 247152 508898 247194 509134
rect 246874 508866 247194 508898
rect 252805 509454 253125 509486
rect 252805 509218 252847 509454
rect 253083 509218 253125 509454
rect 252805 509134 253125 509218
rect 252805 508898 252847 509134
rect 253083 508898 253125 509134
rect 252805 508866 253125 508898
rect 274874 509454 275194 509486
rect 274874 509218 274916 509454
rect 275152 509218 275194 509454
rect 274874 509134 275194 509218
rect 274874 508898 274916 509134
rect 275152 508898 275194 509134
rect 274874 508866 275194 508898
rect 280805 509454 281125 509486
rect 280805 509218 280847 509454
rect 281083 509218 281125 509454
rect 280805 509134 281125 509218
rect 280805 508898 280847 509134
rect 281083 508898 281125 509134
rect 280805 508866 281125 508898
rect 302874 509454 303194 509486
rect 302874 509218 302916 509454
rect 303152 509218 303194 509454
rect 302874 509134 303194 509218
rect 302874 508898 302916 509134
rect 303152 508898 303194 509134
rect 302874 508866 303194 508898
rect 308805 509454 309125 509486
rect 308805 509218 308847 509454
rect 309083 509218 309125 509454
rect 308805 509134 309125 509218
rect 308805 508898 308847 509134
rect 309083 508898 309125 509134
rect 308805 508866 309125 508898
rect 330874 509454 331194 509486
rect 330874 509218 330916 509454
rect 331152 509218 331194 509454
rect 330874 509134 331194 509218
rect 330874 508898 330916 509134
rect 331152 508898 331194 509134
rect 330874 508866 331194 508898
rect 336805 509454 337125 509486
rect 336805 509218 336847 509454
rect 337083 509218 337125 509454
rect 336805 509134 337125 509218
rect 336805 508898 336847 509134
rect 337083 508898 337125 509134
rect 336805 508866 337125 508898
rect 358874 509454 359194 509486
rect 358874 509218 358916 509454
rect 359152 509218 359194 509454
rect 358874 509134 359194 509218
rect 358874 508898 358916 509134
rect 359152 508898 359194 509134
rect 358874 508866 359194 508898
rect 364805 509454 365125 509486
rect 364805 509218 364847 509454
rect 365083 509218 365125 509454
rect 364805 509134 365125 509218
rect 364805 508898 364847 509134
rect 365083 508898 365125 509134
rect 364805 508866 365125 508898
rect 386874 509454 387194 509486
rect 386874 509218 386916 509454
rect 387152 509218 387194 509454
rect 386874 509134 387194 509218
rect 386874 508898 386916 509134
rect 387152 508898 387194 509134
rect 386874 508866 387194 508898
rect 392805 509454 393125 509486
rect 392805 509218 392847 509454
rect 393083 509218 393125 509454
rect 392805 509134 393125 509218
rect 392805 508898 392847 509134
rect 393083 508898 393125 509134
rect 392805 508866 393125 508898
rect 414874 509454 415194 509486
rect 414874 509218 414916 509454
rect 415152 509218 415194 509454
rect 414874 509134 415194 509218
rect 414874 508898 414916 509134
rect 415152 508898 415194 509134
rect 414874 508866 415194 508898
rect 420805 509454 421125 509486
rect 420805 509218 420847 509454
rect 421083 509218 421125 509454
rect 420805 509134 421125 509218
rect 420805 508898 420847 509134
rect 421083 508898 421125 509134
rect 420805 508866 421125 508898
rect 442874 509454 443194 509486
rect 442874 509218 442916 509454
rect 443152 509218 443194 509454
rect 442874 509134 443194 509218
rect 442874 508898 442916 509134
rect 443152 508898 443194 509134
rect 442874 508866 443194 508898
rect 448805 509454 449125 509486
rect 448805 509218 448847 509454
rect 449083 509218 449125 509454
rect 448805 509134 449125 509218
rect 448805 508898 448847 509134
rect 449083 508898 449125 509134
rect 448805 508866 449125 508898
rect 470874 509454 471194 509486
rect 470874 509218 470916 509454
rect 471152 509218 471194 509454
rect 470874 509134 471194 509218
rect 470874 508898 470916 509134
rect 471152 508898 471194 509134
rect 470874 508866 471194 508898
rect 476805 509454 477125 509486
rect 476805 509218 476847 509454
rect 477083 509218 477125 509454
rect 476805 509134 477125 509218
rect 476805 508898 476847 509134
rect 477083 508898 477125 509134
rect 476805 508866 477125 508898
rect 498874 509454 499194 509486
rect 498874 509218 498916 509454
rect 499152 509218 499194 509454
rect 498874 509134 499194 509218
rect 498874 508898 498916 509134
rect 499152 508898 499194 509134
rect 498874 508866 499194 508898
rect 504805 509454 505125 509486
rect 504805 509218 504847 509454
rect 505083 509218 505125 509454
rect 504805 509134 505125 509218
rect 504805 508898 504847 509134
rect 505083 508898 505125 509134
rect 504805 508866 505125 508898
rect 526874 509454 527194 509486
rect 526874 509218 526916 509454
rect 527152 509218 527194 509454
rect 526874 509134 527194 509218
rect 526874 508898 526916 509134
rect 527152 508898 527194 509134
rect 526874 508866 527194 508898
rect 532805 509454 533125 509486
rect 532805 509218 532847 509454
rect 533083 509218 533125 509454
rect 532805 509134 533125 509218
rect 532805 508898 532847 509134
rect 533083 508898 533125 509134
rect 532805 508866 533125 508898
rect 554874 509454 555194 509486
rect 554874 509218 554916 509454
rect 555152 509218 555194 509454
rect 554874 509134 555194 509218
rect 554874 508898 554916 509134
rect 555152 508898 555194 509134
rect 554874 508866 555194 508898
rect 560805 509454 561125 509486
rect 560805 509218 560847 509454
rect 561083 509218 561125 509454
rect 560805 509134 561125 509218
rect 560805 508898 560847 509134
rect 561083 508898 561125 509134
rect 560805 508866 561125 508898
rect -2006 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 -1386 485829
rect -2006 485509 -1386 485593
rect -2006 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 -1386 485509
rect -2006 458829 -1386 485273
rect 19910 485829 20230 485861
rect 19910 485593 19952 485829
rect 20188 485593 20230 485829
rect 19910 485509 20230 485593
rect 19910 485273 19952 485509
rect 20188 485273 20230 485509
rect 19910 485241 20230 485273
rect 25840 485829 26160 485861
rect 25840 485593 25882 485829
rect 26118 485593 26160 485829
rect 25840 485509 26160 485593
rect 25840 485273 25882 485509
rect 26118 485273 26160 485509
rect 25840 485241 26160 485273
rect 31771 485829 32091 485861
rect 31771 485593 31813 485829
rect 32049 485593 32091 485829
rect 31771 485509 32091 485593
rect 31771 485273 31813 485509
rect 32049 485273 32091 485509
rect 31771 485241 32091 485273
rect 47910 485829 48230 485861
rect 47910 485593 47952 485829
rect 48188 485593 48230 485829
rect 47910 485509 48230 485593
rect 47910 485273 47952 485509
rect 48188 485273 48230 485509
rect 47910 485241 48230 485273
rect 53840 485829 54160 485861
rect 53840 485593 53882 485829
rect 54118 485593 54160 485829
rect 53840 485509 54160 485593
rect 53840 485273 53882 485509
rect 54118 485273 54160 485509
rect 53840 485241 54160 485273
rect 59771 485829 60091 485861
rect 59771 485593 59813 485829
rect 60049 485593 60091 485829
rect 59771 485509 60091 485593
rect 59771 485273 59813 485509
rect 60049 485273 60091 485509
rect 59771 485241 60091 485273
rect 75910 485829 76230 485861
rect 75910 485593 75952 485829
rect 76188 485593 76230 485829
rect 75910 485509 76230 485593
rect 75910 485273 75952 485509
rect 76188 485273 76230 485509
rect 75910 485241 76230 485273
rect 81840 485829 82160 485861
rect 81840 485593 81882 485829
rect 82118 485593 82160 485829
rect 81840 485509 82160 485593
rect 81840 485273 81882 485509
rect 82118 485273 82160 485509
rect 81840 485241 82160 485273
rect 87771 485829 88091 485861
rect 87771 485593 87813 485829
rect 88049 485593 88091 485829
rect 87771 485509 88091 485593
rect 87771 485273 87813 485509
rect 88049 485273 88091 485509
rect 87771 485241 88091 485273
rect 103910 485829 104230 485861
rect 103910 485593 103952 485829
rect 104188 485593 104230 485829
rect 103910 485509 104230 485593
rect 103910 485273 103952 485509
rect 104188 485273 104230 485509
rect 103910 485241 104230 485273
rect 109840 485829 110160 485861
rect 109840 485593 109882 485829
rect 110118 485593 110160 485829
rect 109840 485509 110160 485593
rect 109840 485273 109882 485509
rect 110118 485273 110160 485509
rect 109840 485241 110160 485273
rect 115771 485829 116091 485861
rect 115771 485593 115813 485829
rect 116049 485593 116091 485829
rect 115771 485509 116091 485593
rect 115771 485273 115813 485509
rect 116049 485273 116091 485509
rect 115771 485241 116091 485273
rect 131910 485829 132230 485861
rect 131910 485593 131952 485829
rect 132188 485593 132230 485829
rect 131910 485509 132230 485593
rect 131910 485273 131952 485509
rect 132188 485273 132230 485509
rect 131910 485241 132230 485273
rect 137840 485829 138160 485861
rect 137840 485593 137882 485829
rect 138118 485593 138160 485829
rect 137840 485509 138160 485593
rect 137840 485273 137882 485509
rect 138118 485273 138160 485509
rect 137840 485241 138160 485273
rect 143771 485829 144091 485861
rect 143771 485593 143813 485829
rect 144049 485593 144091 485829
rect 143771 485509 144091 485593
rect 143771 485273 143813 485509
rect 144049 485273 144091 485509
rect 143771 485241 144091 485273
rect 159910 485829 160230 485861
rect 159910 485593 159952 485829
rect 160188 485593 160230 485829
rect 159910 485509 160230 485593
rect 159910 485273 159952 485509
rect 160188 485273 160230 485509
rect 159910 485241 160230 485273
rect 165840 485829 166160 485861
rect 165840 485593 165882 485829
rect 166118 485593 166160 485829
rect 165840 485509 166160 485593
rect 165840 485273 165882 485509
rect 166118 485273 166160 485509
rect 165840 485241 166160 485273
rect 171771 485829 172091 485861
rect 171771 485593 171813 485829
rect 172049 485593 172091 485829
rect 171771 485509 172091 485593
rect 171771 485273 171813 485509
rect 172049 485273 172091 485509
rect 171771 485241 172091 485273
rect 187910 485829 188230 485861
rect 187910 485593 187952 485829
rect 188188 485593 188230 485829
rect 187910 485509 188230 485593
rect 187910 485273 187952 485509
rect 188188 485273 188230 485509
rect 187910 485241 188230 485273
rect 193840 485829 194160 485861
rect 193840 485593 193882 485829
rect 194118 485593 194160 485829
rect 193840 485509 194160 485593
rect 193840 485273 193882 485509
rect 194118 485273 194160 485509
rect 193840 485241 194160 485273
rect 199771 485829 200091 485861
rect 199771 485593 199813 485829
rect 200049 485593 200091 485829
rect 199771 485509 200091 485593
rect 199771 485273 199813 485509
rect 200049 485273 200091 485509
rect 199771 485241 200091 485273
rect 215910 485829 216230 485861
rect 215910 485593 215952 485829
rect 216188 485593 216230 485829
rect 215910 485509 216230 485593
rect 215910 485273 215952 485509
rect 216188 485273 216230 485509
rect 215910 485241 216230 485273
rect 221840 485829 222160 485861
rect 221840 485593 221882 485829
rect 222118 485593 222160 485829
rect 221840 485509 222160 485593
rect 221840 485273 221882 485509
rect 222118 485273 222160 485509
rect 221840 485241 222160 485273
rect 227771 485829 228091 485861
rect 227771 485593 227813 485829
rect 228049 485593 228091 485829
rect 227771 485509 228091 485593
rect 227771 485273 227813 485509
rect 228049 485273 228091 485509
rect 227771 485241 228091 485273
rect 243910 485829 244230 485861
rect 243910 485593 243952 485829
rect 244188 485593 244230 485829
rect 243910 485509 244230 485593
rect 243910 485273 243952 485509
rect 244188 485273 244230 485509
rect 243910 485241 244230 485273
rect 249840 485829 250160 485861
rect 249840 485593 249882 485829
rect 250118 485593 250160 485829
rect 249840 485509 250160 485593
rect 249840 485273 249882 485509
rect 250118 485273 250160 485509
rect 249840 485241 250160 485273
rect 255771 485829 256091 485861
rect 255771 485593 255813 485829
rect 256049 485593 256091 485829
rect 255771 485509 256091 485593
rect 255771 485273 255813 485509
rect 256049 485273 256091 485509
rect 255771 485241 256091 485273
rect 271910 485829 272230 485861
rect 271910 485593 271952 485829
rect 272188 485593 272230 485829
rect 271910 485509 272230 485593
rect 271910 485273 271952 485509
rect 272188 485273 272230 485509
rect 271910 485241 272230 485273
rect 277840 485829 278160 485861
rect 277840 485593 277882 485829
rect 278118 485593 278160 485829
rect 277840 485509 278160 485593
rect 277840 485273 277882 485509
rect 278118 485273 278160 485509
rect 277840 485241 278160 485273
rect 283771 485829 284091 485861
rect 283771 485593 283813 485829
rect 284049 485593 284091 485829
rect 283771 485509 284091 485593
rect 283771 485273 283813 485509
rect 284049 485273 284091 485509
rect 283771 485241 284091 485273
rect 299910 485829 300230 485861
rect 299910 485593 299952 485829
rect 300188 485593 300230 485829
rect 299910 485509 300230 485593
rect 299910 485273 299952 485509
rect 300188 485273 300230 485509
rect 299910 485241 300230 485273
rect 305840 485829 306160 485861
rect 305840 485593 305882 485829
rect 306118 485593 306160 485829
rect 305840 485509 306160 485593
rect 305840 485273 305882 485509
rect 306118 485273 306160 485509
rect 305840 485241 306160 485273
rect 311771 485829 312091 485861
rect 311771 485593 311813 485829
rect 312049 485593 312091 485829
rect 311771 485509 312091 485593
rect 311771 485273 311813 485509
rect 312049 485273 312091 485509
rect 311771 485241 312091 485273
rect 327910 485829 328230 485861
rect 327910 485593 327952 485829
rect 328188 485593 328230 485829
rect 327910 485509 328230 485593
rect 327910 485273 327952 485509
rect 328188 485273 328230 485509
rect 327910 485241 328230 485273
rect 333840 485829 334160 485861
rect 333840 485593 333882 485829
rect 334118 485593 334160 485829
rect 333840 485509 334160 485593
rect 333840 485273 333882 485509
rect 334118 485273 334160 485509
rect 333840 485241 334160 485273
rect 339771 485829 340091 485861
rect 339771 485593 339813 485829
rect 340049 485593 340091 485829
rect 339771 485509 340091 485593
rect 339771 485273 339813 485509
rect 340049 485273 340091 485509
rect 339771 485241 340091 485273
rect 355910 485829 356230 485861
rect 355910 485593 355952 485829
rect 356188 485593 356230 485829
rect 355910 485509 356230 485593
rect 355910 485273 355952 485509
rect 356188 485273 356230 485509
rect 355910 485241 356230 485273
rect 361840 485829 362160 485861
rect 361840 485593 361882 485829
rect 362118 485593 362160 485829
rect 361840 485509 362160 485593
rect 361840 485273 361882 485509
rect 362118 485273 362160 485509
rect 361840 485241 362160 485273
rect 367771 485829 368091 485861
rect 367771 485593 367813 485829
rect 368049 485593 368091 485829
rect 367771 485509 368091 485593
rect 367771 485273 367813 485509
rect 368049 485273 368091 485509
rect 367771 485241 368091 485273
rect 383910 485829 384230 485861
rect 383910 485593 383952 485829
rect 384188 485593 384230 485829
rect 383910 485509 384230 485593
rect 383910 485273 383952 485509
rect 384188 485273 384230 485509
rect 383910 485241 384230 485273
rect 389840 485829 390160 485861
rect 389840 485593 389882 485829
rect 390118 485593 390160 485829
rect 389840 485509 390160 485593
rect 389840 485273 389882 485509
rect 390118 485273 390160 485509
rect 389840 485241 390160 485273
rect 395771 485829 396091 485861
rect 395771 485593 395813 485829
rect 396049 485593 396091 485829
rect 395771 485509 396091 485593
rect 395771 485273 395813 485509
rect 396049 485273 396091 485509
rect 395771 485241 396091 485273
rect 411910 485829 412230 485861
rect 411910 485593 411952 485829
rect 412188 485593 412230 485829
rect 411910 485509 412230 485593
rect 411910 485273 411952 485509
rect 412188 485273 412230 485509
rect 411910 485241 412230 485273
rect 417840 485829 418160 485861
rect 417840 485593 417882 485829
rect 418118 485593 418160 485829
rect 417840 485509 418160 485593
rect 417840 485273 417882 485509
rect 418118 485273 418160 485509
rect 417840 485241 418160 485273
rect 423771 485829 424091 485861
rect 423771 485593 423813 485829
rect 424049 485593 424091 485829
rect 423771 485509 424091 485593
rect 423771 485273 423813 485509
rect 424049 485273 424091 485509
rect 423771 485241 424091 485273
rect 439910 485829 440230 485861
rect 439910 485593 439952 485829
rect 440188 485593 440230 485829
rect 439910 485509 440230 485593
rect 439910 485273 439952 485509
rect 440188 485273 440230 485509
rect 439910 485241 440230 485273
rect 445840 485829 446160 485861
rect 445840 485593 445882 485829
rect 446118 485593 446160 485829
rect 445840 485509 446160 485593
rect 445840 485273 445882 485509
rect 446118 485273 446160 485509
rect 445840 485241 446160 485273
rect 451771 485829 452091 485861
rect 451771 485593 451813 485829
rect 452049 485593 452091 485829
rect 451771 485509 452091 485593
rect 451771 485273 451813 485509
rect 452049 485273 452091 485509
rect 451771 485241 452091 485273
rect 467910 485829 468230 485861
rect 467910 485593 467952 485829
rect 468188 485593 468230 485829
rect 467910 485509 468230 485593
rect 467910 485273 467952 485509
rect 468188 485273 468230 485509
rect 467910 485241 468230 485273
rect 473840 485829 474160 485861
rect 473840 485593 473882 485829
rect 474118 485593 474160 485829
rect 473840 485509 474160 485593
rect 473840 485273 473882 485509
rect 474118 485273 474160 485509
rect 473840 485241 474160 485273
rect 479771 485829 480091 485861
rect 479771 485593 479813 485829
rect 480049 485593 480091 485829
rect 479771 485509 480091 485593
rect 479771 485273 479813 485509
rect 480049 485273 480091 485509
rect 479771 485241 480091 485273
rect 495910 485829 496230 485861
rect 495910 485593 495952 485829
rect 496188 485593 496230 485829
rect 495910 485509 496230 485593
rect 495910 485273 495952 485509
rect 496188 485273 496230 485509
rect 495910 485241 496230 485273
rect 501840 485829 502160 485861
rect 501840 485593 501882 485829
rect 502118 485593 502160 485829
rect 501840 485509 502160 485593
rect 501840 485273 501882 485509
rect 502118 485273 502160 485509
rect 501840 485241 502160 485273
rect 507771 485829 508091 485861
rect 507771 485593 507813 485829
rect 508049 485593 508091 485829
rect 507771 485509 508091 485593
rect 507771 485273 507813 485509
rect 508049 485273 508091 485509
rect 507771 485241 508091 485273
rect 523910 485829 524230 485861
rect 523910 485593 523952 485829
rect 524188 485593 524230 485829
rect 523910 485509 524230 485593
rect 523910 485273 523952 485509
rect 524188 485273 524230 485509
rect 523910 485241 524230 485273
rect 529840 485829 530160 485861
rect 529840 485593 529882 485829
rect 530118 485593 530160 485829
rect 529840 485509 530160 485593
rect 529840 485273 529882 485509
rect 530118 485273 530160 485509
rect 529840 485241 530160 485273
rect 535771 485829 536091 485861
rect 535771 485593 535813 485829
rect 536049 485593 536091 485829
rect 535771 485509 536091 485593
rect 535771 485273 535813 485509
rect 536049 485273 536091 485509
rect 535771 485241 536091 485273
rect 551910 485829 552230 485861
rect 551910 485593 551952 485829
rect 552188 485593 552230 485829
rect 551910 485509 552230 485593
rect 551910 485273 551952 485509
rect 552188 485273 552230 485509
rect 551910 485241 552230 485273
rect 557840 485829 558160 485861
rect 557840 485593 557882 485829
rect 558118 485593 558160 485829
rect 557840 485509 558160 485593
rect 557840 485273 557882 485509
rect 558118 485273 558160 485509
rect 557840 485241 558160 485273
rect 563771 485829 564091 485861
rect 563771 485593 563813 485829
rect 564049 485593 564091 485829
rect 563771 485509 564091 485593
rect 563771 485273 563813 485509
rect 564049 485273 564091 485509
rect 563771 485241 564091 485273
rect 573494 485829 574114 512273
rect 573494 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 574114 485829
rect 573494 485509 574114 485593
rect 573494 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 574114 485509
rect 22874 482454 23194 482486
rect 22874 482218 22916 482454
rect 23152 482218 23194 482454
rect 22874 482134 23194 482218
rect 22874 481898 22916 482134
rect 23152 481898 23194 482134
rect 22874 481866 23194 481898
rect 28805 482454 29125 482486
rect 28805 482218 28847 482454
rect 29083 482218 29125 482454
rect 28805 482134 29125 482218
rect 28805 481898 28847 482134
rect 29083 481898 29125 482134
rect 28805 481866 29125 481898
rect 50874 482454 51194 482486
rect 50874 482218 50916 482454
rect 51152 482218 51194 482454
rect 50874 482134 51194 482218
rect 50874 481898 50916 482134
rect 51152 481898 51194 482134
rect 50874 481866 51194 481898
rect 56805 482454 57125 482486
rect 56805 482218 56847 482454
rect 57083 482218 57125 482454
rect 56805 482134 57125 482218
rect 56805 481898 56847 482134
rect 57083 481898 57125 482134
rect 56805 481866 57125 481898
rect 78874 482454 79194 482486
rect 78874 482218 78916 482454
rect 79152 482218 79194 482454
rect 78874 482134 79194 482218
rect 78874 481898 78916 482134
rect 79152 481898 79194 482134
rect 78874 481866 79194 481898
rect 84805 482454 85125 482486
rect 84805 482218 84847 482454
rect 85083 482218 85125 482454
rect 84805 482134 85125 482218
rect 84805 481898 84847 482134
rect 85083 481898 85125 482134
rect 84805 481866 85125 481898
rect 106874 482454 107194 482486
rect 106874 482218 106916 482454
rect 107152 482218 107194 482454
rect 106874 482134 107194 482218
rect 106874 481898 106916 482134
rect 107152 481898 107194 482134
rect 106874 481866 107194 481898
rect 112805 482454 113125 482486
rect 112805 482218 112847 482454
rect 113083 482218 113125 482454
rect 112805 482134 113125 482218
rect 112805 481898 112847 482134
rect 113083 481898 113125 482134
rect 112805 481866 113125 481898
rect 134874 482454 135194 482486
rect 134874 482218 134916 482454
rect 135152 482218 135194 482454
rect 134874 482134 135194 482218
rect 134874 481898 134916 482134
rect 135152 481898 135194 482134
rect 134874 481866 135194 481898
rect 140805 482454 141125 482486
rect 140805 482218 140847 482454
rect 141083 482218 141125 482454
rect 140805 482134 141125 482218
rect 140805 481898 140847 482134
rect 141083 481898 141125 482134
rect 140805 481866 141125 481898
rect 162874 482454 163194 482486
rect 162874 482218 162916 482454
rect 163152 482218 163194 482454
rect 162874 482134 163194 482218
rect 162874 481898 162916 482134
rect 163152 481898 163194 482134
rect 162874 481866 163194 481898
rect 168805 482454 169125 482486
rect 168805 482218 168847 482454
rect 169083 482218 169125 482454
rect 168805 482134 169125 482218
rect 168805 481898 168847 482134
rect 169083 481898 169125 482134
rect 168805 481866 169125 481898
rect 190874 482454 191194 482486
rect 190874 482218 190916 482454
rect 191152 482218 191194 482454
rect 190874 482134 191194 482218
rect 190874 481898 190916 482134
rect 191152 481898 191194 482134
rect 190874 481866 191194 481898
rect 196805 482454 197125 482486
rect 196805 482218 196847 482454
rect 197083 482218 197125 482454
rect 196805 482134 197125 482218
rect 196805 481898 196847 482134
rect 197083 481898 197125 482134
rect 196805 481866 197125 481898
rect 218874 482454 219194 482486
rect 218874 482218 218916 482454
rect 219152 482218 219194 482454
rect 218874 482134 219194 482218
rect 218874 481898 218916 482134
rect 219152 481898 219194 482134
rect 218874 481866 219194 481898
rect 224805 482454 225125 482486
rect 224805 482218 224847 482454
rect 225083 482218 225125 482454
rect 224805 482134 225125 482218
rect 224805 481898 224847 482134
rect 225083 481898 225125 482134
rect 224805 481866 225125 481898
rect 246874 482454 247194 482486
rect 246874 482218 246916 482454
rect 247152 482218 247194 482454
rect 246874 482134 247194 482218
rect 246874 481898 246916 482134
rect 247152 481898 247194 482134
rect 246874 481866 247194 481898
rect 252805 482454 253125 482486
rect 252805 482218 252847 482454
rect 253083 482218 253125 482454
rect 252805 482134 253125 482218
rect 252805 481898 252847 482134
rect 253083 481898 253125 482134
rect 252805 481866 253125 481898
rect 274874 482454 275194 482486
rect 274874 482218 274916 482454
rect 275152 482218 275194 482454
rect 274874 482134 275194 482218
rect 274874 481898 274916 482134
rect 275152 481898 275194 482134
rect 274874 481866 275194 481898
rect 280805 482454 281125 482486
rect 280805 482218 280847 482454
rect 281083 482218 281125 482454
rect 280805 482134 281125 482218
rect 280805 481898 280847 482134
rect 281083 481898 281125 482134
rect 280805 481866 281125 481898
rect 302874 482454 303194 482486
rect 302874 482218 302916 482454
rect 303152 482218 303194 482454
rect 302874 482134 303194 482218
rect 302874 481898 302916 482134
rect 303152 481898 303194 482134
rect 302874 481866 303194 481898
rect 308805 482454 309125 482486
rect 308805 482218 308847 482454
rect 309083 482218 309125 482454
rect 308805 482134 309125 482218
rect 308805 481898 308847 482134
rect 309083 481898 309125 482134
rect 308805 481866 309125 481898
rect 330874 482454 331194 482486
rect 330874 482218 330916 482454
rect 331152 482218 331194 482454
rect 330874 482134 331194 482218
rect 330874 481898 330916 482134
rect 331152 481898 331194 482134
rect 330874 481866 331194 481898
rect 336805 482454 337125 482486
rect 336805 482218 336847 482454
rect 337083 482218 337125 482454
rect 336805 482134 337125 482218
rect 336805 481898 336847 482134
rect 337083 481898 337125 482134
rect 336805 481866 337125 481898
rect 358874 482454 359194 482486
rect 358874 482218 358916 482454
rect 359152 482218 359194 482454
rect 358874 482134 359194 482218
rect 358874 481898 358916 482134
rect 359152 481898 359194 482134
rect 358874 481866 359194 481898
rect 364805 482454 365125 482486
rect 364805 482218 364847 482454
rect 365083 482218 365125 482454
rect 364805 482134 365125 482218
rect 364805 481898 364847 482134
rect 365083 481898 365125 482134
rect 364805 481866 365125 481898
rect 386874 482454 387194 482486
rect 386874 482218 386916 482454
rect 387152 482218 387194 482454
rect 386874 482134 387194 482218
rect 386874 481898 386916 482134
rect 387152 481898 387194 482134
rect 386874 481866 387194 481898
rect 392805 482454 393125 482486
rect 392805 482218 392847 482454
rect 393083 482218 393125 482454
rect 392805 482134 393125 482218
rect 392805 481898 392847 482134
rect 393083 481898 393125 482134
rect 392805 481866 393125 481898
rect 414874 482454 415194 482486
rect 414874 482218 414916 482454
rect 415152 482218 415194 482454
rect 414874 482134 415194 482218
rect 414874 481898 414916 482134
rect 415152 481898 415194 482134
rect 414874 481866 415194 481898
rect 420805 482454 421125 482486
rect 420805 482218 420847 482454
rect 421083 482218 421125 482454
rect 420805 482134 421125 482218
rect 420805 481898 420847 482134
rect 421083 481898 421125 482134
rect 420805 481866 421125 481898
rect 442874 482454 443194 482486
rect 442874 482218 442916 482454
rect 443152 482218 443194 482454
rect 442874 482134 443194 482218
rect 442874 481898 442916 482134
rect 443152 481898 443194 482134
rect 442874 481866 443194 481898
rect 448805 482454 449125 482486
rect 448805 482218 448847 482454
rect 449083 482218 449125 482454
rect 448805 482134 449125 482218
rect 448805 481898 448847 482134
rect 449083 481898 449125 482134
rect 448805 481866 449125 481898
rect 470874 482454 471194 482486
rect 470874 482218 470916 482454
rect 471152 482218 471194 482454
rect 470874 482134 471194 482218
rect 470874 481898 470916 482134
rect 471152 481898 471194 482134
rect 470874 481866 471194 481898
rect 476805 482454 477125 482486
rect 476805 482218 476847 482454
rect 477083 482218 477125 482454
rect 476805 482134 477125 482218
rect 476805 481898 476847 482134
rect 477083 481898 477125 482134
rect 476805 481866 477125 481898
rect 498874 482454 499194 482486
rect 498874 482218 498916 482454
rect 499152 482218 499194 482454
rect 498874 482134 499194 482218
rect 498874 481898 498916 482134
rect 499152 481898 499194 482134
rect 498874 481866 499194 481898
rect 504805 482454 505125 482486
rect 504805 482218 504847 482454
rect 505083 482218 505125 482454
rect 504805 482134 505125 482218
rect 504805 481898 504847 482134
rect 505083 481898 505125 482134
rect 504805 481866 505125 481898
rect 526874 482454 527194 482486
rect 526874 482218 526916 482454
rect 527152 482218 527194 482454
rect 526874 482134 527194 482218
rect 526874 481898 526916 482134
rect 527152 481898 527194 482134
rect 526874 481866 527194 481898
rect 532805 482454 533125 482486
rect 532805 482218 532847 482454
rect 533083 482218 533125 482454
rect 532805 482134 533125 482218
rect 532805 481898 532847 482134
rect 533083 481898 533125 482134
rect 532805 481866 533125 481898
rect 554874 482454 555194 482486
rect 554874 482218 554916 482454
rect 555152 482218 555194 482454
rect 554874 482134 555194 482218
rect 554874 481898 554916 482134
rect 555152 481898 555194 482134
rect 554874 481866 555194 481898
rect 560805 482454 561125 482486
rect 560805 482218 560847 482454
rect 561083 482218 561125 482454
rect 560805 482134 561125 482218
rect 560805 481898 560847 482134
rect 561083 481898 561125 482134
rect 560805 481866 561125 481898
rect -2006 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 -1386 458829
rect -2006 458509 -1386 458593
rect -2006 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 -1386 458509
rect -2006 431829 -1386 458273
rect 19910 458829 20230 458861
rect 19910 458593 19952 458829
rect 20188 458593 20230 458829
rect 19910 458509 20230 458593
rect 19910 458273 19952 458509
rect 20188 458273 20230 458509
rect 19910 458241 20230 458273
rect 25840 458829 26160 458861
rect 25840 458593 25882 458829
rect 26118 458593 26160 458829
rect 25840 458509 26160 458593
rect 25840 458273 25882 458509
rect 26118 458273 26160 458509
rect 25840 458241 26160 458273
rect 31771 458829 32091 458861
rect 31771 458593 31813 458829
rect 32049 458593 32091 458829
rect 31771 458509 32091 458593
rect 31771 458273 31813 458509
rect 32049 458273 32091 458509
rect 31771 458241 32091 458273
rect 47910 458829 48230 458861
rect 47910 458593 47952 458829
rect 48188 458593 48230 458829
rect 47910 458509 48230 458593
rect 47910 458273 47952 458509
rect 48188 458273 48230 458509
rect 47910 458241 48230 458273
rect 53840 458829 54160 458861
rect 53840 458593 53882 458829
rect 54118 458593 54160 458829
rect 53840 458509 54160 458593
rect 53840 458273 53882 458509
rect 54118 458273 54160 458509
rect 53840 458241 54160 458273
rect 59771 458829 60091 458861
rect 59771 458593 59813 458829
rect 60049 458593 60091 458829
rect 59771 458509 60091 458593
rect 59771 458273 59813 458509
rect 60049 458273 60091 458509
rect 59771 458241 60091 458273
rect 75910 458829 76230 458861
rect 75910 458593 75952 458829
rect 76188 458593 76230 458829
rect 75910 458509 76230 458593
rect 75910 458273 75952 458509
rect 76188 458273 76230 458509
rect 75910 458241 76230 458273
rect 81840 458829 82160 458861
rect 81840 458593 81882 458829
rect 82118 458593 82160 458829
rect 81840 458509 82160 458593
rect 81840 458273 81882 458509
rect 82118 458273 82160 458509
rect 81840 458241 82160 458273
rect 87771 458829 88091 458861
rect 87771 458593 87813 458829
rect 88049 458593 88091 458829
rect 87771 458509 88091 458593
rect 87771 458273 87813 458509
rect 88049 458273 88091 458509
rect 87771 458241 88091 458273
rect 103910 458829 104230 458861
rect 103910 458593 103952 458829
rect 104188 458593 104230 458829
rect 103910 458509 104230 458593
rect 103910 458273 103952 458509
rect 104188 458273 104230 458509
rect 103910 458241 104230 458273
rect 109840 458829 110160 458861
rect 109840 458593 109882 458829
rect 110118 458593 110160 458829
rect 109840 458509 110160 458593
rect 109840 458273 109882 458509
rect 110118 458273 110160 458509
rect 109840 458241 110160 458273
rect 115771 458829 116091 458861
rect 115771 458593 115813 458829
rect 116049 458593 116091 458829
rect 115771 458509 116091 458593
rect 115771 458273 115813 458509
rect 116049 458273 116091 458509
rect 115771 458241 116091 458273
rect 131910 458829 132230 458861
rect 131910 458593 131952 458829
rect 132188 458593 132230 458829
rect 131910 458509 132230 458593
rect 131910 458273 131952 458509
rect 132188 458273 132230 458509
rect 131910 458241 132230 458273
rect 137840 458829 138160 458861
rect 137840 458593 137882 458829
rect 138118 458593 138160 458829
rect 137840 458509 138160 458593
rect 137840 458273 137882 458509
rect 138118 458273 138160 458509
rect 137840 458241 138160 458273
rect 143771 458829 144091 458861
rect 143771 458593 143813 458829
rect 144049 458593 144091 458829
rect 143771 458509 144091 458593
rect 143771 458273 143813 458509
rect 144049 458273 144091 458509
rect 143771 458241 144091 458273
rect 159910 458829 160230 458861
rect 159910 458593 159952 458829
rect 160188 458593 160230 458829
rect 159910 458509 160230 458593
rect 159910 458273 159952 458509
rect 160188 458273 160230 458509
rect 159910 458241 160230 458273
rect 165840 458829 166160 458861
rect 165840 458593 165882 458829
rect 166118 458593 166160 458829
rect 165840 458509 166160 458593
rect 165840 458273 165882 458509
rect 166118 458273 166160 458509
rect 165840 458241 166160 458273
rect 171771 458829 172091 458861
rect 171771 458593 171813 458829
rect 172049 458593 172091 458829
rect 171771 458509 172091 458593
rect 171771 458273 171813 458509
rect 172049 458273 172091 458509
rect 171771 458241 172091 458273
rect 187910 458829 188230 458861
rect 187910 458593 187952 458829
rect 188188 458593 188230 458829
rect 187910 458509 188230 458593
rect 187910 458273 187952 458509
rect 188188 458273 188230 458509
rect 187910 458241 188230 458273
rect 193840 458829 194160 458861
rect 193840 458593 193882 458829
rect 194118 458593 194160 458829
rect 193840 458509 194160 458593
rect 193840 458273 193882 458509
rect 194118 458273 194160 458509
rect 193840 458241 194160 458273
rect 199771 458829 200091 458861
rect 199771 458593 199813 458829
rect 200049 458593 200091 458829
rect 199771 458509 200091 458593
rect 199771 458273 199813 458509
rect 200049 458273 200091 458509
rect 199771 458241 200091 458273
rect 215910 458829 216230 458861
rect 215910 458593 215952 458829
rect 216188 458593 216230 458829
rect 215910 458509 216230 458593
rect 215910 458273 215952 458509
rect 216188 458273 216230 458509
rect 215910 458241 216230 458273
rect 221840 458829 222160 458861
rect 221840 458593 221882 458829
rect 222118 458593 222160 458829
rect 221840 458509 222160 458593
rect 221840 458273 221882 458509
rect 222118 458273 222160 458509
rect 221840 458241 222160 458273
rect 227771 458829 228091 458861
rect 227771 458593 227813 458829
rect 228049 458593 228091 458829
rect 227771 458509 228091 458593
rect 227771 458273 227813 458509
rect 228049 458273 228091 458509
rect 227771 458241 228091 458273
rect 243910 458829 244230 458861
rect 243910 458593 243952 458829
rect 244188 458593 244230 458829
rect 243910 458509 244230 458593
rect 243910 458273 243952 458509
rect 244188 458273 244230 458509
rect 243910 458241 244230 458273
rect 249840 458829 250160 458861
rect 249840 458593 249882 458829
rect 250118 458593 250160 458829
rect 249840 458509 250160 458593
rect 249840 458273 249882 458509
rect 250118 458273 250160 458509
rect 249840 458241 250160 458273
rect 255771 458829 256091 458861
rect 255771 458593 255813 458829
rect 256049 458593 256091 458829
rect 255771 458509 256091 458593
rect 255771 458273 255813 458509
rect 256049 458273 256091 458509
rect 255771 458241 256091 458273
rect 271910 458829 272230 458861
rect 271910 458593 271952 458829
rect 272188 458593 272230 458829
rect 271910 458509 272230 458593
rect 271910 458273 271952 458509
rect 272188 458273 272230 458509
rect 271910 458241 272230 458273
rect 277840 458829 278160 458861
rect 277840 458593 277882 458829
rect 278118 458593 278160 458829
rect 277840 458509 278160 458593
rect 277840 458273 277882 458509
rect 278118 458273 278160 458509
rect 277840 458241 278160 458273
rect 283771 458829 284091 458861
rect 283771 458593 283813 458829
rect 284049 458593 284091 458829
rect 283771 458509 284091 458593
rect 283771 458273 283813 458509
rect 284049 458273 284091 458509
rect 283771 458241 284091 458273
rect 299910 458829 300230 458861
rect 299910 458593 299952 458829
rect 300188 458593 300230 458829
rect 299910 458509 300230 458593
rect 299910 458273 299952 458509
rect 300188 458273 300230 458509
rect 299910 458241 300230 458273
rect 305840 458829 306160 458861
rect 305840 458593 305882 458829
rect 306118 458593 306160 458829
rect 305840 458509 306160 458593
rect 305840 458273 305882 458509
rect 306118 458273 306160 458509
rect 305840 458241 306160 458273
rect 311771 458829 312091 458861
rect 311771 458593 311813 458829
rect 312049 458593 312091 458829
rect 311771 458509 312091 458593
rect 311771 458273 311813 458509
rect 312049 458273 312091 458509
rect 311771 458241 312091 458273
rect 327910 458829 328230 458861
rect 327910 458593 327952 458829
rect 328188 458593 328230 458829
rect 327910 458509 328230 458593
rect 327910 458273 327952 458509
rect 328188 458273 328230 458509
rect 327910 458241 328230 458273
rect 333840 458829 334160 458861
rect 333840 458593 333882 458829
rect 334118 458593 334160 458829
rect 333840 458509 334160 458593
rect 333840 458273 333882 458509
rect 334118 458273 334160 458509
rect 333840 458241 334160 458273
rect 339771 458829 340091 458861
rect 339771 458593 339813 458829
rect 340049 458593 340091 458829
rect 339771 458509 340091 458593
rect 339771 458273 339813 458509
rect 340049 458273 340091 458509
rect 339771 458241 340091 458273
rect 355910 458829 356230 458861
rect 355910 458593 355952 458829
rect 356188 458593 356230 458829
rect 355910 458509 356230 458593
rect 355910 458273 355952 458509
rect 356188 458273 356230 458509
rect 355910 458241 356230 458273
rect 361840 458829 362160 458861
rect 361840 458593 361882 458829
rect 362118 458593 362160 458829
rect 361840 458509 362160 458593
rect 361840 458273 361882 458509
rect 362118 458273 362160 458509
rect 361840 458241 362160 458273
rect 367771 458829 368091 458861
rect 367771 458593 367813 458829
rect 368049 458593 368091 458829
rect 367771 458509 368091 458593
rect 367771 458273 367813 458509
rect 368049 458273 368091 458509
rect 367771 458241 368091 458273
rect 383910 458829 384230 458861
rect 383910 458593 383952 458829
rect 384188 458593 384230 458829
rect 383910 458509 384230 458593
rect 383910 458273 383952 458509
rect 384188 458273 384230 458509
rect 383910 458241 384230 458273
rect 389840 458829 390160 458861
rect 389840 458593 389882 458829
rect 390118 458593 390160 458829
rect 389840 458509 390160 458593
rect 389840 458273 389882 458509
rect 390118 458273 390160 458509
rect 389840 458241 390160 458273
rect 395771 458829 396091 458861
rect 395771 458593 395813 458829
rect 396049 458593 396091 458829
rect 395771 458509 396091 458593
rect 395771 458273 395813 458509
rect 396049 458273 396091 458509
rect 395771 458241 396091 458273
rect 411910 458829 412230 458861
rect 411910 458593 411952 458829
rect 412188 458593 412230 458829
rect 411910 458509 412230 458593
rect 411910 458273 411952 458509
rect 412188 458273 412230 458509
rect 411910 458241 412230 458273
rect 417840 458829 418160 458861
rect 417840 458593 417882 458829
rect 418118 458593 418160 458829
rect 417840 458509 418160 458593
rect 417840 458273 417882 458509
rect 418118 458273 418160 458509
rect 417840 458241 418160 458273
rect 423771 458829 424091 458861
rect 423771 458593 423813 458829
rect 424049 458593 424091 458829
rect 423771 458509 424091 458593
rect 423771 458273 423813 458509
rect 424049 458273 424091 458509
rect 423771 458241 424091 458273
rect 439910 458829 440230 458861
rect 439910 458593 439952 458829
rect 440188 458593 440230 458829
rect 439910 458509 440230 458593
rect 439910 458273 439952 458509
rect 440188 458273 440230 458509
rect 439910 458241 440230 458273
rect 445840 458829 446160 458861
rect 445840 458593 445882 458829
rect 446118 458593 446160 458829
rect 445840 458509 446160 458593
rect 445840 458273 445882 458509
rect 446118 458273 446160 458509
rect 445840 458241 446160 458273
rect 451771 458829 452091 458861
rect 451771 458593 451813 458829
rect 452049 458593 452091 458829
rect 451771 458509 452091 458593
rect 451771 458273 451813 458509
rect 452049 458273 452091 458509
rect 451771 458241 452091 458273
rect 467910 458829 468230 458861
rect 467910 458593 467952 458829
rect 468188 458593 468230 458829
rect 467910 458509 468230 458593
rect 467910 458273 467952 458509
rect 468188 458273 468230 458509
rect 467910 458241 468230 458273
rect 473840 458829 474160 458861
rect 473840 458593 473882 458829
rect 474118 458593 474160 458829
rect 473840 458509 474160 458593
rect 473840 458273 473882 458509
rect 474118 458273 474160 458509
rect 473840 458241 474160 458273
rect 479771 458829 480091 458861
rect 479771 458593 479813 458829
rect 480049 458593 480091 458829
rect 479771 458509 480091 458593
rect 479771 458273 479813 458509
rect 480049 458273 480091 458509
rect 479771 458241 480091 458273
rect 495910 458829 496230 458861
rect 495910 458593 495952 458829
rect 496188 458593 496230 458829
rect 495910 458509 496230 458593
rect 495910 458273 495952 458509
rect 496188 458273 496230 458509
rect 495910 458241 496230 458273
rect 501840 458829 502160 458861
rect 501840 458593 501882 458829
rect 502118 458593 502160 458829
rect 501840 458509 502160 458593
rect 501840 458273 501882 458509
rect 502118 458273 502160 458509
rect 501840 458241 502160 458273
rect 507771 458829 508091 458861
rect 507771 458593 507813 458829
rect 508049 458593 508091 458829
rect 507771 458509 508091 458593
rect 507771 458273 507813 458509
rect 508049 458273 508091 458509
rect 507771 458241 508091 458273
rect 523910 458829 524230 458861
rect 523910 458593 523952 458829
rect 524188 458593 524230 458829
rect 523910 458509 524230 458593
rect 523910 458273 523952 458509
rect 524188 458273 524230 458509
rect 523910 458241 524230 458273
rect 529840 458829 530160 458861
rect 529840 458593 529882 458829
rect 530118 458593 530160 458829
rect 529840 458509 530160 458593
rect 529840 458273 529882 458509
rect 530118 458273 530160 458509
rect 529840 458241 530160 458273
rect 535771 458829 536091 458861
rect 535771 458593 535813 458829
rect 536049 458593 536091 458829
rect 535771 458509 536091 458593
rect 535771 458273 535813 458509
rect 536049 458273 536091 458509
rect 535771 458241 536091 458273
rect 551910 458829 552230 458861
rect 551910 458593 551952 458829
rect 552188 458593 552230 458829
rect 551910 458509 552230 458593
rect 551910 458273 551952 458509
rect 552188 458273 552230 458509
rect 551910 458241 552230 458273
rect 557840 458829 558160 458861
rect 557840 458593 557882 458829
rect 558118 458593 558160 458829
rect 557840 458509 558160 458593
rect 557840 458273 557882 458509
rect 558118 458273 558160 458509
rect 557840 458241 558160 458273
rect 563771 458829 564091 458861
rect 563771 458593 563813 458829
rect 564049 458593 564091 458829
rect 563771 458509 564091 458593
rect 563771 458273 563813 458509
rect 564049 458273 564091 458509
rect 563771 458241 564091 458273
rect 573494 458829 574114 485273
rect 573494 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 574114 458829
rect 573494 458509 574114 458593
rect 573494 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 574114 458509
rect 22874 455454 23194 455486
rect 22874 455218 22916 455454
rect 23152 455218 23194 455454
rect 22874 455134 23194 455218
rect 22874 454898 22916 455134
rect 23152 454898 23194 455134
rect 22874 454866 23194 454898
rect 28805 455454 29125 455486
rect 28805 455218 28847 455454
rect 29083 455218 29125 455454
rect 28805 455134 29125 455218
rect 28805 454898 28847 455134
rect 29083 454898 29125 455134
rect 28805 454866 29125 454898
rect 50874 455454 51194 455486
rect 50874 455218 50916 455454
rect 51152 455218 51194 455454
rect 50874 455134 51194 455218
rect 50874 454898 50916 455134
rect 51152 454898 51194 455134
rect 50874 454866 51194 454898
rect 56805 455454 57125 455486
rect 56805 455218 56847 455454
rect 57083 455218 57125 455454
rect 56805 455134 57125 455218
rect 56805 454898 56847 455134
rect 57083 454898 57125 455134
rect 56805 454866 57125 454898
rect 78874 455454 79194 455486
rect 78874 455218 78916 455454
rect 79152 455218 79194 455454
rect 78874 455134 79194 455218
rect 78874 454898 78916 455134
rect 79152 454898 79194 455134
rect 78874 454866 79194 454898
rect 84805 455454 85125 455486
rect 84805 455218 84847 455454
rect 85083 455218 85125 455454
rect 84805 455134 85125 455218
rect 84805 454898 84847 455134
rect 85083 454898 85125 455134
rect 84805 454866 85125 454898
rect 106874 455454 107194 455486
rect 106874 455218 106916 455454
rect 107152 455218 107194 455454
rect 106874 455134 107194 455218
rect 106874 454898 106916 455134
rect 107152 454898 107194 455134
rect 106874 454866 107194 454898
rect 112805 455454 113125 455486
rect 112805 455218 112847 455454
rect 113083 455218 113125 455454
rect 112805 455134 113125 455218
rect 112805 454898 112847 455134
rect 113083 454898 113125 455134
rect 112805 454866 113125 454898
rect 134874 455454 135194 455486
rect 134874 455218 134916 455454
rect 135152 455218 135194 455454
rect 134874 455134 135194 455218
rect 134874 454898 134916 455134
rect 135152 454898 135194 455134
rect 134874 454866 135194 454898
rect 140805 455454 141125 455486
rect 140805 455218 140847 455454
rect 141083 455218 141125 455454
rect 140805 455134 141125 455218
rect 140805 454898 140847 455134
rect 141083 454898 141125 455134
rect 140805 454866 141125 454898
rect 162874 455454 163194 455486
rect 162874 455218 162916 455454
rect 163152 455218 163194 455454
rect 162874 455134 163194 455218
rect 162874 454898 162916 455134
rect 163152 454898 163194 455134
rect 162874 454866 163194 454898
rect 168805 455454 169125 455486
rect 168805 455218 168847 455454
rect 169083 455218 169125 455454
rect 168805 455134 169125 455218
rect 168805 454898 168847 455134
rect 169083 454898 169125 455134
rect 168805 454866 169125 454898
rect 190874 455454 191194 455486
rect 190874 455218 190916 455454
rect 191152 455218 191194 455454
rect 190874 455134 191194 455218
rect 190874 454898 190916 455134
rect 191152 454898 191194 455134
rect 190874 454866 191194 454898
rect 196805 455454 197125 455486
rect 196805 455218 196847 455454
rect 197083 455218 197125 455454
rect 196805 455134 197125 455218
rect 196805 454898 196847 455134
rect 197083 454898 197125 455134
rect 196805 454866 197125 454898
rect 218874 455454 219194 455486
rect 218874 455218 218916 455454
rect 219152 455218 219194 455454
rect 218874 455134 219194 455218
rect 218874 454898 218916 455134
rect 219152 454898 219194 455134
rect 218874 454866 219194 454898
rect 224805 455454 225125 455486
rect 224805 455218 224847 455454
rect 225083 455218 225125 455454
rect 224805 455134 225125 455218
rect 224805 454898 224847 455134
rect 225083 454898 225125 455134
rect 224805 454866 225125 454898
rect 246874 455454 247194 455486
rect 246874 455218 246916 455454
rect 247152 455218 247194 455454
rect 246874 455134 247194 455218
rect 246874 454898 246916 455134
rect 247152 454898 247194 455134
rect 246874 454866 247194 454898
rect 252805 455454 253125 455486
rect 252805 455218 252847 455454
rect 253083 455218 253125 455454
rect 252805 455134 253125 455218
rect 252805 454898 252847 455134
rect 253083 454898 253125 455134
rect 252805 454866 253125 454898
rect 274874 455454 275194 455486
rect 274874 455218 274916 455454
rect 275152 455218 275194 455454
rect 274874 455134 275194 455218
rect 274874 454898 274916 455134
rect 275152 454898 275194 455134
rect 274874 454866 275194 454898
rect 280805 455454 281125 455486
rect 280805 455218 280847 455454
rect 281083 455218 281125 455454
rect 280805 455134 281125 455218
rect 280805 454898 280847 455134
rect 281083 454898 281125 455134
rect 280805 454866 281125 454898
rect 302874 455454 303194 455486
rect 302874 455218 302916 455454
rect 303152 455218 303194 455454
rect 302874 455134 303194 455218
rect 302874 454898 302916 455134
rect 303152 454898 303194 455134
rect 302874 454866 303194 454898
rect 308805 455454 309125 455486
rect 308805 455218 308847 455454
rect 309083 455218 309125 455454
rect 308805 455134 309125 455218
rect 308805 454898 308847 455134
rect 309083 454898 309125 455134
rect 308805 454866 309125 454898
rect 330874 455454 331194 455486
rect 330874 455218 330916 455454
rect 331152 455218 331194 455454
rect 330874 455134 331194 455218
rect 330874 454898 330916 455134
rect 331152 454898 331194 455134
rect 330874 454866 331194 454898
rect 336805 455454 337125 455486
rect 336805 455218 336847 455454
rect 337083 455218 337125 455454
rect 336805 455134 337125 455218
rect 336805 454898 336847 455134
rect 337083 454898 337125 455134
rect 336805 454866 337125 454898
rect 358874 455454 359194 455486
rect 358874 455218 358916 455454
rect 359152 455218 359194 455454
rect 358874 455134 359194 455218
rect 358874 454898 358916 455134
rect 359152 454898 359194 455134
rect 358874 454866 359194 454898
rect 364805 455454 365125 455486
rect 364805 455218 364847 455454
rect 365083 455218 365125 455454
rect 364805 455134 365125 455218
rect 364805 454898 364847 455134
rect 365083 454898 365125 455134
rect 364805 454866 365125 454898
rect 386874 455454 387194 455486
rect 386874 455218 386916 455454
rect 387152 455218 387194 455454
rect 386874 455134 387194 455218
rect 386874 454898 386916 455134
rect 387152 454898 387194 455134
rect 386874 454866 387194 454898
rect 392805 455454 393125 455486
rect 392805 455218 392847 455454
rect 393083 455218 393125 455454
rect 392805 455134 393125 455218
rect 392805 454898 392847 455134
rect 393083 454898 393125 455134
rect 392805 454866 393125 454898
rect 414874 455454 415194 455486
rect 414874 455218 414916 455454
rect 415152 455218 415194 455454
rect 414874 455134 415194 455218
rect 414874 454898 414916 455134
rect 415152 454898 415194 455134
rect 414874 454866 415194 454898
rect 420805 455454 421125 455486
rect 420805 455218 420847 455454
rect 421083 455218 421125 455454
rect 420805 455134 421125 455218
rect 420805 454898 420847 455134
rect 421083 454898 421125 455134
rect 420805 454866 421125 454898
rect 442874 455454 443194 455486
rect 442874 455218 442916 455454
rect 443152 455218 443194 455454
rect 442874 455134 443194 455218
rect 442874 454898 442916 455134
rect 443152 454898 443194 455134
rect 442874 454866 443194 454898
rect 448805 455454 449125 455486
rect 448805 455218 448847 455454
rect 449083 455218 449125 455454
rect 448805 455134 449125 455218
rect 448805 454898 448847 455134
rect 449083 454898 449125 455134
rect 448805 454866 449125 454898
rect 470874 455454 471194 455486
rect 470874 455218 470916 455454
rect 471152 455218 471194 455454
rect 470874 455134 471194 455218
rect 470874 454898 470916 455134
rect 471152 454898 471194 455134
rect 470874 454866 471194 454898
rect 476805 455454 477125 455486
rect 476805 455218 476847 455454
rect 477083 455218 477125 455454
rect 476805 455134 477125 455218
rect 476805 454898 476847 455134
rect 477083 454898 477125 455134
rect 476805 454866 477125 454898
rect 498874 455454 499194 455486
rect 498874 455218 498916 455454
rect 499152 455218 499194 455454
rect 498874 455134 499194 455218
rect 498874 454898 498916 455134
rect 499152 454898 499194 455134
rect 498874 454866 499194 454898
rect 504805 455454 505125 455486
rect 504805 455218 504847 455454
rect 505083 455218 505125 455454
rect 504805 455134 505125 455218
rect 504805 454898 504847 455134
rect 505083 454898 505125 455134
rect 504805 454866 505125 454898
rect 526874 455454 527194 455486
rect 526874 455218 526916 455454
rect 527152 455218 527194 455454
rect 526874 455134 527194 455218
rect 526874 454898 526916 455134
rect 527152 454898 527194 455134
rect 526874 454866 527194 454898
rect 532805 455454 533125 455486
rect 532805 455218 532847 455454
rect 533083 455218 533125 455454
rect 532805 455134 533125 455218
rect 532805 454898 532847 455134
rect 533083 454898 533125 455134
rect 532805 454866 533125 454898
rect 554874 455454 555194 455486
rect 554874 455218 554916 455454
rect 555152 455218 555194 455454
rect 554874 455134 555194 455218
rect 554874 454898 554916 455134
rect 555152 454898 555194 455134
rect 554874 454866 555194 454898
rect 560805 455454 561125 455486
rect 560805 455218 560847 455454
rect 561083 455218 561125 455454
rect 560805 455134 561125 455218
rect 560805 454898 560847 455134
rect 561083 454898 561125 455134
rect 560805 454866 561125 454898
rect -2006 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 -1386 431829
rect -2006 431509 -1386 431593
rect -2006 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 -1386 431509
rect -2006 404829 -1386 431273
rect 19910 431829 20230 431861
rect 19910 431593 19952 431829
rect 20188 431593 20230 431829
rect 19910 431509 20230 431593
rect 19910 431273 19952 431509
rect 20188 431273 20230 431509
rect 19910 431241 20230 431273
rect 25840 431829 26160 431861
rect 25840 431593 25882 431829
rect 26118 431593 26160 431829
rect 25840 431509 26160 431593
rect 25840 431273 25882 431509
rect 26118 431273 26160 431509
rect 25840 431241 26160 431273
rect 31771 431829 32091 431861
rect 31771 431593 31813 431829
rect 32049 431593 32091 431829
rect 31771 431509 32091 431593
rect 31771 431273 31813 431509
rect 32049 431273 32091 431509
rect 31771 431241 32091 431273
rect 47910 431829 48230 431861
rect 47910 431593 47952 431829
rect 48188 431593 48230 431829
rect 47910 431509 48230 431593
rect 47910 431273 47952 431509
rect 48188 431273 48230 431509
rect 47910 431241 48230 431273
rect 53840 431829 54160 431861
rect 53840 431593 53882 431829
rect 54118 431593 54160 431829
rect 53840 431509 54160 431593
rect 53840 431273 53882 431509
rect 54118 431273 54160 431509
rect 53840 431241 54160 431273
rect 59771 431829 60091 431861
rect 59771 431593 59813 431829
rect 60049 431593 60091 431829
rect 59771 431509 60091 431593
rect 59771 431273 59813 431509
rect 60049 431273 60091 431509
rect 59771 431241 60091 431273
rect 75910 431829 76230 431861
rect 75910 431593 75952 431829
rect 76188 431593 76230 431829
rect 75910 431509 76230 431593
rect 75910 431273 75952 431509
rect 76188 431273 76230 431509
rect 75910 431241 76230 431273
rect 81840 431829 82160 431861
rect 81840 431593 81882 431829
rect 82118 431593 82160 431829
rect 81840 431509 82160 431593
rect 81840 431273 81882 431509
rect 82118 431273 82160 431509
rect 81840 431241 82160 431273
rect 87771 431829 88091 431861
rect 87771 431593 87813 431829
rect 88049 431593 88091 431829
rect 87771 431509 88091 431593
rect 87771 431273 87813 431509
rect 88049 431273 88091 431509
rect 87771 431241 88091 431273
rect 103910 431829 104230 431861
rect 103910 431593 103952 431829
rect 104188 431593 104230 431829
rect 103910 431509 104230 431593
rect 103910 431273 103952 431509
rect 104188 431273 104230 431509
rect 103910 431241 104230 431273
rect 109840 431829 110160 431861
rect 109840 431593 109882 431829
rect 110118 431593 110160 431829
rect 109840 431509 110160 431593
rect 109840 431273 109882 431509
rect 110118 431273 110160 431509
rect 109840 431241 110160 431273
rect 115771 431829 116091 431861
rect 115771 431593 115813 431829
rect 116049 431593 116091 431829
rect 115771 431509 116091 431593
rect 115771 431273 115813 431509
rect 116049 431273 116091 431509
rect 115771 431241 116091 431273
rect 131910 431829 132230 431861
rect 131910 431593 131952 431829
rect 132188 431593 132230 431829
rect 131910 431509 132230 431593
rect 131910 431273 131952 431509
rect 132188 431273 132230 431509
rect 131910 431241 132230 431273
rect 137840 431829 138160 431861
rect 137840 431593 137882 431829
rect 138118 431593 138160 431829
rect 137840 431509 138160 431593
rect 137840 431273 137882 431509
rect 138118 431273 138160 431509
rect 137840 431241 138160 431273
rect 143771 431829 144091 431861
rect 143771 431593 143813 431829
rect 144049 431593 144091 431829
rect 143771 431509 144091 431593
rect 143771 431273 143813 431509
rect 144049 431273 144091 431509
rect 143771 431241 144091 431273
rect 159910 431829 160230 431861
rect 159910 431593 159952 431829
rect 160188 431593 160230 431829
rect 159910 431509 160230 431593
rect 159910 431273 159952 431509
rect 160188 431273 160230 431509
rect 159910 431241 160230 431273
rect 165840 431829 166160 431861
rect 165840 431593 165882 431829
rect 166118 431593 166160 431829
rect 165840 431509 166160 431593
rect 165840 431273 165882 431509
rect 166118 431273 166160 431509
rect 165840 431241 166160 431273
rect 171771 431829 172091 431861
rect 171771 431593 171813 431829
rect 172049 431593 172091 431829
rect 171771 431509 172091 431593
rect 171771 431273 171813 431509
rect 172049 431273 172091 431509
rect 171771 431241 172091 431273
rect 187910 431829 188230 431861
rect 187910 431593 187952 431829
rect 188188 431593 188230 431829
rect 187910 431509 188230 431593
rect 187910 431273 187952 431509
rect 188188 431273 188230 431509
rect 187910 431241 188230 431273
rect 193840 431829 194160 431861
rect 193840 431593 193882 431829
rect 194118 431593 194160 431829
rect 193840 431509 194160 431593
rect 193840 431273 193882 431509
rect 194118 431273 194160 431509
rect 193840 431241 194160 431273
rect 199771 431829 200091 431861
rect 199771 431593 199813 431829
rect 200049 431593 200091 431829
rect 199771 431509 200091 431593
rect 199771 431273 199813 431509
rect 200049 431273 200091 431509
rect 199771 431241 200091 431273
rect 215910 431829 216230 431861
rect 215910 431593 215952 431829
rect 216188 431593 216230 431829
rect 215910 431509 216230 431593
rect 215910 431273 215952 431509
rect 216188 431273 216230 431509
rect 215910 431241 216230 431273
rect 221840 431829 222160 431861
rect 221840 431593 221882 431829
rect 222118 431593 222160 431829
rect 221840 431509 222160 431593
rect 221840 431273 221882 431509
rect 222118 431273 222160 431509
rect 221840 431241 222160 431273
rect 227771 431829 228091 431861
rect 227771 431593 227813 431829
rect 228049 431593 228091 431829
rect 227771 431509 228091 431593
rect 227771 431273 227813 431509
rect 228049 431273 228091 431509
rect 227771 431241 228091 431273
rect 243910 431829 244230 431861
rect 243910 431593 243952 431829
rect 244188 431593 244230 431829
rect 243910 431509 244230 431593
rect 243910 431273 243952 431509
rect 244188 431273 244230 431509
rect 243910 431241 244230 431273
rect 249840 431829 250160 431861
rect 249840 431593 249882 431829
rect 250118 431593 250160 431829
rect 249840 431509 250160 431593
rect 249840 431273 249882 431509
rect 250118 431273 250160 431509
rect 249840 431241 250160 431273
rect 255771 431829 256091 431861
rect 255771 431593 255813 431829
rect 256049 431593 256091 431829
rect 255771 431509 256091 431593
rect 255771 431273 255813 431509
rect 256049 431273 256091 431509
rect 255771 431241 256091 431273
rect 271910 431829 272230 431861
rect 271910 431593 271952 431829
rect 272188 431593 272230 431829
rect 271910 431509 272230 431593
rect 271910 431273 271952 431509
rect 272188 431273 272230 431509
rect 271910 431241 272230 431273
rect 277840 431829 278160 431861
rect 277840 431593 277882 431829
rect 278118 431593 278160 431829
rect 277840 431509 278160 431593
rect 277840 431273 277882 431509
rect 278118 431273 278160 431509
rect 277840 431241 278160 431273
rect 283771 431829 284091 431861
rect 283771 431593 283813 431829
rect 284049 431593 284091 431829
rect 283771 431509 284091 431593
rect 283771 431273 283813 431509
rect 284049 431273 284091 431509
rect 283771 431241 284091 431273
rect 299910 431829 300230 431861
rect 299910 431593 299952 431829
rect 300188 431593 300230 431829
rect 299910 431509 300230 431593
rect 299910 431273 299952 431509
rect 300188 431273 300230 431509
rect 299910 431241 300230 431273
rect 305840 431829 306160 431861
rect 305840 431593 305882 431829
rect 306118 431593 306160 431829
rect 305840 431509 306160 431593
rect 305840 431273 305882 431509
rect 306118 431273 306160 431509
rect 305840 431241 306160 431273
rect 311771 431829 312091 431861
rect 311771 431593 311813 431829
rect 312049 431593 312091 431829
rect 311771 431509 312091 431593
rect 311771 431273 311813 431509
rect 312049 431273 312091 431509
rect 311771 431241 312091 431273
rect 327910 431829 328230 431861
rect 327910 431593 327952 431829
rect 328188 431593 328230 431829
rect 327910 431509 328230 431593
rect 327910 431273 327952 431509
rect 328188 431273 328230 431509
rect 327910 431241 328230 431273
rect 333840 431829 334160 431861
rect 333840 431593 333882 431829
rect 334118 431593 334160 431829
rect 333840 431509 334160 431593
rect 333840 431273 333882 431509
rect 334118 431273 334160 431509
rect 333840 431241 334160 431273
rect 339771 431829 340091 431861
rect 339771 431593 339813 431829
rect 340049 431593 340091 431829
rect 339771 431509 340091 431593
rect 339771 431273 339813 431509
rect 340049 431273 340091 431509
rect 339771 431241 340091 431273
rect 355910 431829 356230 431861
rect 355910 431593 355952 431829
rect 356188 431593 356230 431829
rect 355910 431509 356230 431593
rect 355910 431273 355952 431509
rect 356188 431273 356230 431509
rect 355910 431241 356230 431273
rect 361840 431829 362160 431861
rect 361840 431593 361882 431829
rect 362118 431593 362160 431829
rect 361840 431509 362160 431593
rect 361840 431273 361882 431509
rect 362118 431273 362160 431509
rect 361840 431241 362160 431273
rect 367771 431829 368091 431861
rect 367771 431593 367813 431829
rect 368049 431593 368091 431829
rect 367771 431509 368091 431593
rect 367771 431273 367813 431509
rect 368049 431273 368091 431509
rect 367771 431241 368091 431273
rect 383910 431829 384230 431861
rect 383910 431593 383952 431829
rect 384188 431593 384230 431829
rect 383910 431509 384230 431593
rect 383910 431273 383952 431509
rect 384188 431273 384230 431509
rect 383910 431241 384230 431273
rect 389840 431829 390160 431861
rect 389840 431593 389882 431829
rect 390118 431593 390160 431829
rect 389840 431509 390160 431593
rect 389840 431273 389882 431509
rect 390118 431273 390160 431509
rect 389840 431241 390160 431273
rect 395771 431829 396091 431861
rect 395771 431593 395813 431829
rect 396049 431593 396091 431829
rect 395771 431509 396091 431593
rect 395771 431273 395813 431509
rect 396049 431273 396091 431509
rect 395771 431241 396091 431273
rect 411910 431829 412230 431861
rect 411910 431593 411952 431829
rect 412188 431593 412230 431829
rect 411910 431509 412230 431593
rect 411910 431273 411952 431509
rect 412188 431273 412230 431509
rect 411910 431241 412230 431273
rect 417840 431829 418160 431861
rect 417840 431593 417882 431829
rect 418118 431593 418160 431829
rect 417840 431509 418160 431593
rect 417840 431273 417882 431509
rect 418118 431273 418160 431509
rect 417840 431241 418160 431273
rect 423771 431829 424091 431861
rect 423771 431593 423813 431829
rect 424049 431593 424091 431829
rect 423771 431509 424091 431593
rect 423771 431273 423813 431509
rect 424049 431273 424091 431509
rect 423771 431241 424091 431273
rect 439910 431829 440230 431861
rect 439910 431593 439952 431829
rect 440188 431593 440230 431829
rect 439910 431509 440230 431593
rect 439910 431273 439952 431509
rect 440188 431273 440230 431509
rect 439910 431241 440230 431273
rect 445840 431829 446160 431861
rect 445840 431593 445882 431829
rect 446118 431593 446160 431829
rect 445840 431509 446160 431593
rect 445840 431273 445882 431509
rect 446118 431273 446160 431509
rect 445840 431241 446160 431273
rect 451771 431829 452091 431861
rect 451771 431593 451813 431829
rect 452049 431593 452091 431829
rect 451771 431509 452091 431593
rect 451771 431273 451813 431509
rect 452049 431273 452091 431509
rect 451771 431241 452091 431273
rect 467910 431829 468230 431861
rect 467910 431593 467952 431829
rect 468188 431593 468230 431829
rect 467910 431509 468230 431593
rect 467910 431273 467952 431509
rect 468188 431273 468230 431509
rect 467910 431241 468230 431273
rect 473840 431829 474160 431861
rect 473840 431593 473882 431829
rect 474118 431593 474160 431829
rect 473840 431509 474160 431593
rect 473840 431273 473882 431509
rect 474118 431273 474160 431509
rect 473840 431241 474160 431273
rect 479771 431829 480091 431861
rect 479771 431593 479813 431829
rect 480049 431593 480091 431829
rect 479771 431509 480091 431593
rect 479771 431273 479813 431509
rect 480049 431273 480091 431509
rect 479771 431241 480091 431273
rect 495910 431829 496230 431861
rect 495910 431593 495952 431829
rect 496188 431593 496230 431829
rect 495910 431509 496230 431593
rect 495910 431273 495952 431509
rect 496188 431273 496230 431509
rect 495910 431241 496230 431273
rect 501840 431829 502160 431861
rect 501840 431593 501882 431829
rect 502118 431593 502160 431829
rect 501840 431509 502160 431593
rect 501840 431273 501882 431509
rect 502118 431273 502160 431509
rect 501840 431241 502160 431273
rect 507771 431829 508091 431861
rect 507771 431593 507813 431829
rect 508049 431593 508091 431829
rect 507771 431509 508091 431593
rect 507771 431273 507813 431509
rect 508049 431273 508091 431509
rect 507771 431241 508091 431273
rect 523910 431829 524230 431861
rect 523910 431593 523952 431829
rect 524188 431593 524230 431829
rect 523910 431509 524230 431593
rect 523910 431273 523952 431509
rect 524188 431273 524230 431509
rect 523910 431241 524230 431273
rect 529840 431829 530160 431861
rect 529840 431593 529882 431829
rect 530118 431593 530160 431829
rect 529840 431509 530160 431593
rect 529840 431273 529882 431509
rect 530118 431273 530160 431509
rect 529840 431241 530160 431273
rect 535771 431829 536091 431861
rect 535771 431593 535813 431829
rect 536049 431593 536091 431829
rect 535771 431509 536091 431593
rect 535771 431273 535813 431509
rect 536049 431273 536091 431509
rect 535771 431241 536091 431273
rect 551910 431829 552230 431861
rect 551910 431593 551952 431829
rect 552188 431593 552230 431829
rect 551910 431509 552230 431593
rect 551910 431273 551952 431509
rect 552188 431273 552230 431509
rect 551910 431241 552230 431273
rect 557840 431829 558160 431861
rect 557840 431593 557882 431829
rect 558118 431593 558160 431829
rect 557840 431509 558160 431593
rect 557840 431273 557882 431509
rect 558118 431273 558160 431509
rect 557840 431241 558160 431273
rect 563771 431829 564091 431861
rect 563771 431593 563813 431829
rect 564049 431593 564091 431829
rect 563771 431509 564091 431593
rect 563771 431273 563813 431509
rect 564049 431273 564091 431509
rect 563771 431241 564091 431273
rect 573494 431829 574114 458273
rect 573494 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 574114 431829
rect 573494 431509 574114 431593
rect 573494 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 574114 431509
rect 22874 428454 23194 428486
rect 22874 428218 22916 428454
rect 23152 428218 23194 428454
rect 22874 428134 23194 428218
rect 22874 427898 22916 428134
rect 23152 427898 23194 428134
rect 22874 427866 23194 427898
rect 28805 428454 29125 428486
rect 28805 428218 28847 428454
rect 29083 428218 29125 428454
rect 28805 428134 29125 428218
rect 28805 427898 28847 428134
rect 29083 427898 29125 428134
rect 28805 427866 29125 427898
rect 50874 428454 51194 428486
rect 50874 428218 50916 428454
rect 51152 428218 51194 428454
rect 50874 428134 51194 428218
rect 50874 427898 50916 428134
rect 51152 427898 51194 428134
rect 50874 427866 51194 427898
rect 56805 428454 57125 428486
rect 56805 428218 56847 428454
rect 57083 428218 57125 428454
rect 56805 428134 57125 428218
rect 56805 427898 56847 428134
rect 57083 427898 57125 428134
rect 56805 427866 57125 427898
rect 78874 428454 79194 428486
rect 78874 428218 78916 428454
rect 79152 428218 79194 428454
rect 78874 428134 79194 428218
rect 78874 427898 78916 428134
rect 79152 427898 79194 428134
rect 78874 427866 79194 427898
rect 84805 428454 85125 428486
rect 84805 428218 84847 428454
rect 85083 428218 85125 428454
rect 84805 428134 85125 428218
rect 84805 427898 84847 428134
rect 85083 427898 85125 428134
rect 84805 427866 85125 427898
rect 106874 428454 107194 428486
rect 106874 428218 106916 428454
rect 107152 428218 107194 428454
rect 106874 428134 107194 428218
rect 106874 427898 106916 428134
rect 107152 427898 107194 428134
rect 106874 427866 107194 427898
rect 112805 428454 113125 428486
rect 112805 428218 112847 428454
rect 113083 428218 113125 428454
rect 112805 428134 113125 428218
rect 112805 427898 112847 428134
rect 113083 427898 113125 428134
rect 112805 427866 113125 427898
rect 134874 428454 135194 428486
rect 134874 428218 134916 428454
rect 135152 428218 135194 428454
rect 134874 428134 135194 428218
rect 134874 427898 134916 428134
rect 135152 427898 135194 428134
rect 134874 427866 135194 427898
rect 140805 428454 141125 428486
rect 140805 428218 140847 428454
rect 141083 428218 141125 428454
rect 140805 428134 141125 428218
rect 140805 427898 140847 428134
rect 141083 427898 141125 428134
rect 140805 427866 141125 427898
rect 162874 428454 163194 428486
rect 162874 428218 162916 428454
rect 163152 428218 163194 428454
rect 162874 428134 163194 428218
rect 162874 427898 162916 428134
rect 163152 427898 163194 428134
rect 162874 427866 163194 427898
rect 168805 428454 169125 428486
rect 168805 428218 168847 428454
rect 169083 428218 169125 428454
rect 168805 428134 169125 428218
rect 168805 427898 168847 428134
rect 169083 427898 169125 428134
rect 168805 427866 169125 427898
rect 190874 428454 191194 428486
rect 190874 428218 190916 428454
rect 191152 428218 191194 428454
rect 190874 428134 191194 428218
rect 190874 427898 190916 428134
rect 191152 427898 191194 428134
rect 190874 427866 191194 427898
rect 196805 428454 197125 428486
rect 196805 428218 196847 428454
rect 197083 428218 197125 428454
rect 196805 428134 197125 428218
rect 196805 427898 196847 428134
rect 197083 427898 197125 428134
rect 196805 427866 197125 427898
rect 218874 428454 219194 428486
rect 218874 428218 218916 428454
rect 219152 428218 219194 428454
rect 218874 428134 219194 428218
rect 218874 427898 218916 428134
rect 219152 427898 219194 428134
rect 218874 427866 219194 427898
rect 224805 428454 225125 428486
rect 224805 428218 224847 428454
rect 225083 428218 225125 428454
rect 224805 428134 225125 428218
rect 224805 427898 224847 428134
rect 225083 427898 225125 428134
rect 224805 427866 225125 427898
rect 246874 428454 247194 428486
rect 246874 428218 246916 428454
rect 247152 428218 247194 428454
rect 246874 428134 247194 428218
rect 246874 427898 246916 428134
rect 247152 427898 247194 428134
rect 246874 427866 247194 427898
rect 252805 428454 253125 428486
rect 252805 428218 252847 428454
rect 253083 428218 253125 428454
rect 252805 428134 253125 428218
rect 252805 427898 252847 428134
rect 253083 427898 253125 428134
rect 252805 427866 253125 427898
rect 274874 428454 275194 428486
rect 274874 428218 274916 428454
rect 275152 428218 275194 428454
rect 274874 428134 275194 428218
rect 274874 427898 274916 428134
rect 275152 427898 275194 428134
rect 274874 427866 275194 427898
rect 280805 428454 281125 428486
rect 280805 428218 280847 428454
rect 281083 428218 281125 428454
rect 280805 428134 281125 428218
rect 280805 427898 280847 428134
rect 281083 427898 281125 428134
rect 280805 427866 281125 427898
rect 302874 428454 303194 428486
rect 302874 428218 302916 428454
rect 303152 428218 303194 428454
rect 302874 428134 303194 428218
rect 302874 427898 302916 428134
rect 303152 427898 303194 428134
rect 302874 427866 303194 427898
rect 308805 428454 309125 428486
rect 308805 428218 308847 428454
rect 309083 428218 309125 428454
rect 308805 428134 309125 428218
rect 308805 427898 308847 428134
rect 309083 427898 309125 428134
rect 308805 427866 309125 427898
rect 330874 428454 331194 428486
rect 330874 428218 330916 428454
rect 331152 428218 331194 428454
rect 330874 428134 331194 428218
rect 330874 427898 330916 428134
rect 331152 427898 331194 428134
rect 330874 427866 331194 427898
rect 336805 428454 337125 428486
rect 336805 428218 336847 428454
rect 337083 428218 337125 428454
rect 336805 428134 337125 428218
rect 336805 427898 336847 428134
rect 337083 427898 337125 428134
rect 336805 427866 337125 427898
rect 358874 428454 359194 428486
rect 358874 428218 358916 428454
rect 359152 428218 359194 428454
rect 358874 428134 359194 428218
rect 358874 427898 358916 428134
rect 359152 427898 359194 428134
rect 358874 427866 359194 427898
rect 364805 428454 365125 428486
rect 364805 428218 364847 428454
rect 365083 428218 365125 428454
rect 364805 428134 365125 428218
rect 364805 427898 364847 428134
rect 365083 427898 365125 428134
rect 364805 427866 365125 427898
rect 386874 428454 387194 428486
rect 386874 428218 386916 428454
rect 387152 428218 387194 428454
rect 386874 428134 387194 428218
rect 386874 427898 386916 428134
rect 387152 427898 387194 428134
rect 386874 427866 387194 427898
rect 392805 428454 393125 428486
rect 392805 428218 392847 428454
rect 393083 428218 393125 428454
rect 392805 428134 393125 428218
rect 392805 427898 392847 428134
rect 393083 427898 393125 428134
rect 392805 427866 393125 427898
rect 414874 428454 415194 428486
rect 414874 428218 414916 428454
rect 415152 428218 415194 428454
rect 414874 428134 415194 428218
rect 414874 427898 414916 428134
rect 415152 427898 415194 428134
rect 414874 427866 415194 427898
rect 420805 428454 421125 428486
rect 420805 428218 420847 428454
rect 421083 428218 421125 428454
rect 420805 428134 421125 428218
rect 420805 427898 420847 428134
rect 421083 427898 421125 428134
rect 420805 427866 421125 427898
rect 442874 428454 443194 428486
rect 442874 428218 442916 428454
rect 443152 428218 443194 428454
rect 442874 428134 443194 428218
rect 442874 427898 442916 428134
rect 443152 427898 443194 428134
rect 442874 427866 443194 427898
rect 448805 428454 449125 428486
rect 448805 428218 448847 428454
rect 449083 428218 449125 428454
rect 448805 428134 449125 428218
rect 448805 427898 448847 428134
rect 449083 427898 449125 428134
rect 448805 427866 449125 427898
rect 470874 428454 471194 428486
rect 470874 428218 470916 428454
rect 471152 428218 471194 428454
rect 470874 428134 471194 428218
rect 470874 427898 470916 428134
rect 471152 427898 471194 428134
rect 470874 427866 471194 427898
rect 476805 428454 477125 428486
rect 476805 428218 476847 428454
rect 477083 428218 477125 428454
rect 476805 428134 477125 428218
rect 476805 427898 476847 428134
rect 477083 427898 477125 428134
rect 476805 427866 477125 427898
rect 498874 428454 499194 428486
rect 498874 428218 498916 428454
rect 499152 428218 499194 428454
rect 498874 428134 499194 428218
rect 498874 427898 498916 428134
rect 499152 427898 499194 428134
rect 498874 427866 499194 427898
rect 504805 428454 505125 428486
rect 504805 428218 504847 428454
rect 505083 428218 505125 428454
rect 504805 428134 505125 428218
rect 504805 427898 504847 428134
rect 505083 427898 505125 428134
rect 504805 427866 505125 427898
rect 526874 428454 527194 428486
rect 526874 428218 526916 428454
rect 527152 428218 527194 428454
rect 526874 428134 527194 428218
rect 526874 427898 526916 428134
rect 527152 427898 527194 428134
rect 526874 427866 527194 427898
rect 532805 428454 533125 428486
rect 532805 428218 532847 428454
rect 533083 428218 533125 428454
rect 532805 428134 533125 428218
rect 532805 427898 532847 428134
rect 533083 427898 533125 428134
rect 532805 427866 533125 427898
rect 554874 428454 555194 428486
rect 554874 428218 554916 428454
rect 555152 428218 555194 428454
rect 554874 428134 555194 428218
rect 554874 427898 554916 428134
rect 555152 427898 555194 428134
rect 554874 427866 555194 427898
rect 560805 428454 561125 428486
rect 560805 428218 560847 428454
rect 561083 428218 561125 428454
rect 560805 428134 561125 428218
rect 560805 427898 560847 428134
rect 561083 427898 561125 428134
rect 560805 427866 561125 427898
rect -2006 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 -1386 404829
rect -2006 404509 -1386 404593
rect -2006 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 -1386 404509
rect -2006 377829 -1386 404273
rect 19910 404829 20230 404861
rect 19910 404593 19952 404829
rect 20188 404593 20230 404829
rect 19910 404509 20230 404593
rect 19910 404273 19952 404509
rect 20188 404273 20230 404509
rect 19910 404241 20230 404273
rect 25840 404829 26160 404861
rect 25840 404593 25882 404829
rect 26118 404593 26160 404829
rect 25840 404509 26160 404593
rect 25840 404273 25882 404509
rect 26118 404273 26160 404509
rect 25840 404241 26160 404273
rect 31771 404829 32091 404861
rect 31771 404593 31813 404829
rect 32049 404593 32091 404829
rect 31771 404509 32091 404593
rect 31771 404273 31813 404509
rect 32049 404273 32091 404509
rect 31771 404241 32091 404273
rect 47910 404829 48230 404861
rect 47910 404593 47952 404829
rect 48188 404593 48230 404829
rect 47910 404509 48230 404593
rect 47910 404273 47952 404509
rect 48188 404273 48230 404509
rect 47910 404241 48230 404273
rect 53840 404829 54160 404861
rect 53840 404593 53882 404829
rect 54118 404593 54160 404829
rect 53840 404509 54160 404593
rect 53840 404273 53882 404509
rect 54118 404273 54160 404509
rect 53840 404241 54160 404273
rect 59771 404829 60091 404861
rect 59771 404593 59813 404829
rect 60049 404593 60091 404829
rect 59771 404509 60091 404593
rect 59771 404273 59813 404509
rect 60049 404273 60091 404509
rect 59771 404241 60091 404273
rect 75910 404829 76230 404861
rect 75910 404593 75952 404829
rect 76188 404593 76230 404829
rect 75910 404509 76230 404593
rect 75910 404273 75952 404509
rect 76188 404273 76230 404509
rect 75910 404241 76230 404273
rect 81840 404829 82160 404861
rect 81840 404593 81882 404829
rect 82118 404593 82160 404829
rect 81840 404509 82160 404593
rect 81840 404273 81882 404509
rect 82118 404273 82160 404509
rect 81840 404241 82160 404273
rect 87771 404829 88091 404861
rect 87771 404593 87813 404829
rect 88049 404593 88091 404829
rect 87771 404509 88091 404593
rect 87771 404273 87813 404509
rect 88049 404273 88091 404509
rect 87771 404241 88091 404273
rect 103910 404829 104230 404861
rect 103910 404593 103952 404829
rect 104188 404593 104230 404829
rect 103910 404509 104230 404593
rect 103910 404273 103952 404509
rect 104188 404273 104230 404509
rect 103910 404241 104230 404273
rect 109840 404829 110160 404861
rect 109840 404593 109882 404829
rect 110118 404593 110160 404829
rect 109840 404509 110160 404593
rect 109840 404273 109882 404509
rect 110118 404273 110160 404509
rect 109840 404241 110160 404273
rect 115771 404829 116091 404861
rect 115771 404593 115813 404829
rect 116049 404593 116091 404829
rect 115771 404509 116091 404593
rect 115771 404273 115813 404509
rect 116049 404273 116091 404509
rect 115771 404241 116091 404273
rect 131910 404829 132230 404861
rect 131910 404593 131952 404829
rect 132188 404593 132230 404829
rect 131910 404509 132230 404593
rect 131910 404273 131952 404509
rect 132188 404273 132230 404509
rect 131910 404241 132230 404273
rect 137840 404829 138160 404861
rect 137840 404593 137882 404829
rect 138118 404593 138160 404829
rect 137840 404509 138160 404593
rect 137840 404273 137882 404509
rect 138118 404273 138160 404509
rect 137840 404241 138160 404273
rect 143771 404829 144091 404861
rect 143771 404593 143813 404829
rect 144049 404593 144091 404829
rect 143771 404509 144091 404593
rect 143771 404273 143813 404509
rect 144049 404273 144091 404509
rect 143771 404241 144091 404273
rect 159910 404829 160230 404861
rect 159910 404593 159952 404829
rect 160188 404593 160230 404829
rect 159910 404509 160230 404593
rect 159910 404273 159952 404509
rect 160188 404273 160230 404509
rect 159910 404241 160230 404273
rect 165840 404829 166160 404861
rect 165840 404593 165882 404829
rect 166118 404593 166160 404829
rect 165840 404509 166160 404593
rect 165840 404273 165882 404509
rect 166118 404273 166160 404509
rect 165840 404241 166160 404273
rect 171771 404829 172091 404861
rect 171771 404593 171813 404829
rect 172049 404593 172091 404829
rect 171771 404509 172091 404593
rect 171771 404273 171813 404509
rect 172049 404273 172091 404509
rect 171771 404241 172091 404273
rect 187910 404829 188230 404861
rect 187910 404593 187952 404829
rect 188188 404593 188230 404829
rect 187910 404509 188230 404593
rect 187910 404273 187952 404509
rect 188188 404273 188230 404509
rect 187910 404241 188230 404273
rect 193840 404829 194160 404861
rect 193840 404593 193882 404829
rect 194118 404593 194160 404829
rect 193840 404509 194160 404593
rect 193840 404273 193882 404509
rect 194118 404273 194160 404509
rect 193840 404241 194160 404273
rect 199771 404829 200091 404861
rect 199771 404593 199813 404829
rect 200049 404593 200091 404829
rect 199771 404509 200091 404593
rect 199771 404273 199813 404509
rect 200049 404273 200091 404509
rect 199771 404241 200091 404273
rect 215910 404829 216230 404861
rect 215910 404593 215952 404829
rect 216188 404593 216230 404829
rect 215910 404509 216230 404593
rect 215910 404273 215952 404509
rect 216188 404273 216230 404509
rect 215910 404241 216230 404273
rect 221840 404829 222160 404861
rect 221840 404593 221882 404829
rect 222118 404593 222160 404829
rect 221840 404509 222160 404593
rect 221840 404273 221882 404509
rect 222118 404273 222160 404509
rect 221840 404241 222160 404273
rect 227771 404829 228091 404861
rect 227771 404593 227813 404829
rect 228049 404593 228091 404829
rect 227771 404509 228091 404593
rect 227771 404273 227813 404509
rect 228049 404273 228091 404509
rect 227771 404241 228091 404273
rect 243910 404829 244230 404861
rect 243910 404593 243952 404829
rect 244188 404593 244230 404829
rect 243910 404509 244230 404593
rect 243910 404273 243952 404509
rect 244188 404273 244230 404509
rect 243910 404241 244230 404273
rect 249840 404829 250160 404861
rect 249840 404593 249882 404829
rect 250118 404593 250160 404829
rect 249840 404509 250160 404593
rect 249840 404273 249882 404509
rect 250118 404273 250160 404509
rect 249840 404241 250160 404273
rect 255771 404829 256091 404861
rect 255771 404593 255813 404829
rect 256049 404593 256091 404829
rect 255771 404509 256091 404593
rect 255771 404273 255813 404509
rect 256049 404273 256091 404509
rect 255771 404241 256091 404273
rect 271910 404829 272230 404861
rect 271910 404593 271952 404829
rect 272188 404593 272230 404829
rect 271910 404509 272230 404593
rect 271910 404273 271952 404509
rect 272188 404273 272230 404509
rect 271910 404241 272230 404273
rect 277840 404829 278160 404861
rect 277840 404593 277882 404829
rect 278118 404593 278160 404829
rect 277840 404509 278160 404593
rect 277840 404273 277882 404509
rect 278118 404273 278160 404509
rect 277840 404241 278160 404273
rect 283771 404829 284091 404861
rect 283771 404593 283813 404829
rect 284049 404593 284091 404829
rect 283771 404509 284091 404593
rect 283771 404273 283813 404509
rect 284049 404273 284091 404509
rect 283771 404241 284091 404273
rect 299910 404829 300230 404861
rect 299910 404593 299952 404829
rect 300188 404593 300230 404829
rect 299910 404509 300230 404593
rect 299910 404273 299952 404509
rect 300188 404273 300230 404509
rect 299910 404241 300230 404273
rect 305840 404829 306160 404861
rect 305840 404593 305882 404829
rect 306118 404593 306160 404829
rect 305840 404509 306160 404593
rect 305840 404273 305882 404509
rect 306118 404273 306160 404509
rect 305840 404241 306160 404273
rect 311771 404829 312091 404861
rect 311771 404593 311813 404829
rect 312049 404593 312091 404829
rect 311771 404509 312091 404593
rect 311771 404273 311813 404509
rect 312049 404273 312091 404509
rect 311771 404241 312091 404273
rect 327910 404829 328230 404861
rect 327910 404593 327952 404829
rect 328188 404593 328230 404829
rect 327910 404509 328230 404593
rect 327910 404273 327952 404509
rect 328188 404273 328230 404509
rect 327910 404241 328230 404273
rect 333840 404829 334160 404861
rect 333840 404593 333882 404829
rect 334118 404593 334160 404829
rect 333840 404509 334160 404593
rect 333840 404273 333882 404509
rect 334118 404273 334160 404509
rect 333840 404241 334160 404273
rect 339771 404829 340091 404861
rect 339771 404593 339813 404829
rect 340049 404593 340091 404829
rect 339771 404509 340091 404593
rect 339771 404273 339813 404509
rect 340049 404273 340091 404509
rect 339771 404241 340091 404273
rect 355910 404829 356230 404861
rect 355910 404593 355952 404829
rect 356188 404593 356230 404829
rect 355910 404509 356230 404593
rect 355910 404273 355952 404509
rect 356188 404273 356230 404509
rect 355910 404241 356230 404273
rect 361840 404829 362160 404861
rect 361840 404593 361882 404829
rect 362118 404593 362160 404829
rect 361840 404509 362160 404593
rect 361840 404273 361882 404509
rect 362118 404273 362160 404509
rect 361840 404241 362160 404273
rect 367771 404829 368091 404861
rect 367771 404593 367813 404829
rect 368049 404593 368091 404829
rect 367771 404509 368091 404593
rect 367771 404273 367813 404509
rect 368049 404273 368091 404509
rect 367771 404241 368091 404273
rect 383910 404829 384230 404861
rect 383910 404593 383952 404829
rect 384188 404593 384230 404829
rect 383910 404509 384230 404593
rect 383910 404273 383952 404509
rect 384188 404273 384230 404509
rect 383910 404241 384230 404273
rect 389840 404829 390160 404861
rect 389840 404593 389882 404829
rect 390118 404593 390160 404829
rect 389840 404509 390160 404593
rect 389840 404273 389882 404509
rect 390118 404273 390160 404509
rect 389840 404241 390160 404273
rect 395771 404829 396091 404861
rect 395771 404593 395813 404829
rect 396049 404593 396091 404829
rect 395771 404509 396091 404593
rect 395771 404273 395813 404509
rect 396049 404273 396091 404509
rect 395771 404241 396091 404273
rect 411910 404829 412230 404861
rect 411910 404593 411952 404829
rect 412188 404593 412230 404829
rect 411910 404509 412230 404593
rect 411910 404273 411952 404509
rect 412188 404273 412230 404509
rect 411910 404241 412230 404273
rect 417840 404829 418160 404861
rect 417840 404593 417882 404829
rect 418118 404593 418160 404829
rect 417840 404509 418160 404593
rect 417840 404273 417882 404509
rect 418118 404273 418160 404509
rect 417840 404241 418160 404273
rect 423771 404829 424091 404861
rect 423771 404593 423813 404829
rect 424049 404593 424091 404829
rect 423771 404509 424091 404593
rect 423771 404273 423813 404509
rect 424049 404273 424091 404509
rect 423771 404241 424091 404273
rect 439910 404829 440230 404861
rect 439910 404593 439952 404829
rect 440188 404593 440230 404829
rect 439910 404509 440230 404593
rect 439910 404273 439952 404509
rect 440188 404273 440230 404509
rect 439910 404241 440230 404273
rect 445840 404829 446160 404861
rect 445840 404593 445882 404829
rect 446118 404593 446160 404829
rect 445840 404509 446160 404593
rect 445840 404273 445882 404509
rect 446118 404273 446160 404509
rect 445840 404241 446160 404273
rect 451771 404829 452091 404861
rect 451771 404593 451813 404829
rect 452049 404593 452091 404829
rect 451771 404509 452091 404593
rect 451771 404273 451813 404509
rect 452049 404273 452091 404509
rect 451771 404241 452091 404273
rect 467910 404829 468230 404861
rect 467910 404593 467952 404829
rect 468188 404593 468230 404829
rect 467910 404509 468230 404593
rect 467910 404273 467952 404509
rect 468188 404273 468230 404509
rect 467910 404241 468230 404273
rect 473840 404829 474160 404861
rect 473840 404593 473882 404829
rect 474118 404593 474160 404829
rect 473840 404509 474160 404593
rect 473840 404273 473882 404509
rect 474118 404273 474160 404509
rect 473840 404241 474160 404273
rect 479771 404829 480091 404861
rect 479771 404593 479813 404829
rect 480049 404593 480091 404829
rect 479771 404509 480091 404593
rect 479771 404273 479813 404509
rect 480049 404273 480091 404509
rect 479771 404241 480091 404273
rect 495910 404829 496230 404861
rect 495910 404593 495952 404829
rect 496188 404593 496230 404829
rect 495910 404509 496230 404593
rect 495910 404273 495952 404509
rect 496188 404273 496230 404509
rect 495910 404241 496230 404273
rect 501840 404829 502160 404861
rect 501840 404593 501882 404829
rect 502118 404593 502160 404829
rect 501840 404509 502160 404593
rect 501840 404273 501882 404509
rect 502118 404273 502160 404509
rect 501840 404241 502160 404273
rect 507771 404829 508091 404861
rect 507771 404593 507813 404829
rect 508049 404593 508091 404829
rect 507771 404509 508091 404593
rect 507771 404273 507813 404509
rect 508049 404273 508091 404509
rect 507771 404241 508091 404273
rect 523910 404829 524230 404861
rect 523910 404593 523952 404829
rect 524188 404593 524230 404829
rect 523910 404509 524230 404593
rect 523910 404273 523952 404509
rect 524188 404273 524230 404509
rect 523910 404241 524230 404273
rect 529840 404829 530160 404861
rect 529840 404593 529882 404829
rect 530118 404593 530160 404829
rect 529840 404509 530160 404593
rect 529840 404273 529882 404509
rect 530118 404273 530160 404509
rect 529840 404241 530160 404273
rect 535771 404829 536091 404861
rect 535771 404593 535813 404829
rect 536049 404593 536091 404829
rect 535771 404509 536091 404593
rect 535771 404273 535813 404509
rect 536049 404273 536091 404509
rect 535771 404241 536091 404273
rect 551910 404829 552230 404861
rect 551910 404593 551952 404829
rect 552188 404593 552230 404829
rect 551910 404509 552230 404593
rect 551910 404273 551952 404509
rect 552188 404273 552230 404509
rect 551910 404241 552230 404273
rect 557840 404829 558160 404861
rect 557840 404593 557882 404829
rect 558118 404593 558160 404829
rect 557840 404509 558160 404593
rect 557840 404273 557882 404509
rect 558118 404273 558160 404509
rect 557840 404241 558160 404273
rect 563771 404829 564091 404861
rect 563771 404593 563813 404829
rect 564049 404593 564091 404829
rect 563771 404509 564091 404593
rect 563771 404273 563813 404509
rect 564049 404273 564091 404509
rect 563771 404241 564091 404273
rect 573494 404829 574114 431273
rect 573494 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 574114 404829
rect 573494 404509 574114 404593
rect 573494 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 574114 404509
rect 22874 401454 23194 401486
rect 22874 401218 22916 401454
rect 23152 401218 23194 401454
rect 22874 401134 23194 401218
rect 22874 400898 22916 401134
rect 23152 400898 23194 401134
rect 22874 400866 23194 400898
rect 28805 401454 29125 401486
rect 28805 401218 28847 401454
rect 29083 401218 29125 401454
rect 28805 401134 29125 401218
rect 28805 400898 28847 401134
rect 29083 400898 29125 401134
rect 28805 400866 29125 400898
rect 50874 401454 51194 401486
rect 50874 401218 50916 401454
rect 51152 401218 51194 401454
rect 50874 401134 51194 401218
rect 50874 400898 50916 401134
rect 51152 400898 51194 401134
rect 50874 400866 51194 400898
rect 56805 401454 57125 401486
rect 56805 401218 56847 401454
rect 57083 401218 57125 401454
rect 56805 401134 57125 401218
rect 56805 400898 56847 401134
rect 57083 400898 57125 401134
rect 56805 400866 57125 400898
rect 78874 401454 79194 401486
rect 78874 401218 78916 401454
rect 79152 401218 79194 401454
rect 78874 401134 79194 401218
rect 78874 400898 78916 401134
rect 79152 400898 79194 401134
rect 78874 400866 79194 400898
rect 84805 401454 85125 401486
rect 84805 401218 84847 401454
rect 85083 401218 85125 401454
rect 84805 401134 85125 401218
rect 84805 400898 84847 401134
rect 85083 400898 85125 401134
rect 84805 400866 85125 400898
rect 106874 401454 107194 401486
rect 106874 401218 106916 401454
rect 107152 401218 107194 401454
rect 106874 401134 107194 401218
rect 106874 400898 106916 401134
rect 107152 400898 107194 401134
rect 106874 400866 107194 400898
rect 112805 401454 113125 401486
rect 112805 401218 112847 401454
rect 113083 401218 113125 401454
rect 112805 401134 113125 401218
rect 112805 400898 112847 401134
rect 113083 400898 113125 401134
rect 112805 400866 113125 400898
rect 134874 401454 135194 401486
rect 134874 401218 134916 401454
rect 135152 401218 135194 401454
rect 134874 401134 135194 401218
rect 134874 400898 134916 401134
rect 135152 400898 135194 401134
rect 134874 400866 135194 400898
rect 140805 401454 141125 401486
rect 140805 401218 140847 401454
rect 141083 401218 141125 401454
rect 140805 401134 141125 401218
rect 140805 400898 140847 401134
rect 141083 400898 141125 401134
rect 140805 400866 141125 400898
rect 162874 401454 163194 401486
rect 162874 401218 162916 401454
rect 163152 401218 163194 401454
rect 162874 401134 163194 401218
rect 162874 400898 162916 401134
rect 163152 400898 163194 401134
rect 162874 400866 163194 400898
rect 168805 401454 169125 401486
rect 168805 401218 168847 401454
rect 169083 401218 169125 401454
rect 168805 401134 169125 401218
rect 168805 400898 168847 401134
rect 169083 400898 169125 401134
rect 168805 400866 169125 400898
rect 190874 401454 191194 401486
rect 190874 401218 190916 401454
rect 191152 401218 191194 401454
rect 190874 401134 191194 401218
rect 190874 400898 190916 401134
rect 191152 400898 191194 401134
rect 190874 400866 191194 400898
rect 196805 401454 197125 401486
rect 196805 401218 196847 401454
rect 197083 401218 197125 401454
rect 196805 401134 197125 401218
rect 196805 400898 196847 401134
rect 197083 400898 197125 401134
rect 196805 400866 197125 400898
rect 218874 401454 219194 401486
rect 218874 401218 218916 401454
rect 219152 401218 219194 401454
rect 218874 401134 219194 401218
rect 218874 400898 218916 401134
rect 219152 400898 219194 401134
rect 218874 400866 219194 400898
rect 224805 401454 225125 401486
rect 224805 401218 224847 401454
rect 225083 401218 225125 401454
rect 224805 401134 225125 401218
rect 224805 400898 224847 401134
rect 225083 400898 225125 401134
rect 224805 400866 225125 400898
rect 246874 401454 247194 401486
rect 246874 401218 246916 401454
rect 247152 401218 247194 401454
rect 246874 401134 247194 401218
rect 246874 400898 246916 401134
rect 247152 400898 247194 401134
rect 246874 400866 247194 400898
rect 252805 401454 253125 401486
rect 252805 401218 252847 401454
rect 253083 401218 253125 401454
rect 252805 401134 253125 401218
rect 252805 400898 252847 401134
rect 253083 400898 253125 401134
rect 252805 400866 253125 400898
rect 274874 401454 275194 401486
rect 274874 401218 274916 401454
rect 275152 401218 275194 401454
rect 274874 401134 275194 401218
rect 274874 400898 274916 401134
rect 275152 400898 275194 401134
rect 274874 400866 275194 400898
rect 280805 401454 281125 401486
rect 280805 401218 280847 401454
rect 281083 401218 281125 401454
rect 280805 401134 281125 401218
rect 280805 400898 280847 401134
rect 281083 400898 281125 401134
rect 280805 400866 281125 400898
rect 302874 401454 303194 401486
rect 302874 401218 302916 401454
rect 303152 401218 303194 401454
rect 302874 401134 303194 401218
rect 302874 400898 302916 401134
rect 303152 400898 303194 401134
rect 302874 400866 303194 400898
rect 308805 401454 309125 401486
rect 308805 401218 308847 401454
rect 309083 401218 309125 401454
rect 308805 401134 309125 401218
rect 308805 400898 308847 401134
rect 309083 400898 309125 401134
rect 308805 400866 309125 400898
rect 330874 401454 331194 401486
rect 330874 401218 330916 401454
rect 331152 401218 331194 401454
rect 330874 401134 331194 401218
rect 330874 400898 330916 401134
rect 331152 400898 331194 401134
rect 330874 400866 331194 400898
rect 336805 401454 337125 401486
rect 336805 401218 336847 401454
rect 337083 401218 337125 401454
rect 336805 401134 337125 401218
rect 336805 400898 336847 401134
rect 337083 400898 337125 401134
rect 336805 400866 337125 400898
rect 358874 401454 359194 401486
rect 358874 401218 358916 401454
rect 359152 401218 359194 401454
rect 358874 401134 359194 401218
rect 358874 400898 358916 401134
rect 359152 400898 359194 401134
rect 358874 400866 359194 400898
rect 364805 401454 365125 401486
rect 364805 401218 364847 401454
rect 365083 401218 365125 401454
rect 364805 401134 365125 401218
rect 364805 400898 364847 401134
rect 365083 400898 365125 401134
rect 364805 400866 365125 400898
rect 386874 401454 387194 401486
rect 386874 401218 386916 401454
rect 387152 401218 387194 401454
rect 386874 401134 387194 401218
rect 386874 400898 386916 401134
rect 387152 400898 387194 401134
rect 386874 400866 387194 400898
rect 392805 401454 393125 401486
rect 392805 401218 392847 401454
rect 393083 401218 393125 401454
rect 392805 401134 393125 401218
rect 392805 400898 392847 401134
rect 393083 400898 393125 401134
rect 392805 400866 393125 400898
rect 414874 401454 415194 401486
rect 414874 401218 414916 401454
rect 415152 401218 415194 401454
rect 414874 401134 415194 401218
rect 414874 400898 414916 401134
rect 415152 400898 415194 401134
rect 414874 400866 415194 400898
rect 420805 401454 421125 401486
rect 420805 401218 420847 401454
rect 421083 401218 421125 401454
rect 420805 401134 421125 401218
rect 420805 400898 420847 401134
rect 421083 400898 421125 401134
rect 420805 400866 421125 400898
rect 442874 401454 443194 401486
rect 442874 401218 442916 401454
rect 443152 401218 443194 401454
rect 442874 401134 443194 401218
rect 442874 400898 442916 401134
rect 443152 400898 443194 401134
rect 442874 400866 443194 400898
rect 448805 401454 449125 401486
rect 448805 401218 448847 401454
rect 449083 401218 449125 401454
rect 448805 401134 449125 401218
rect 448805 400898 448847 401134
rect 449083 400898 449125 401134
rect 448805 400866 449125 400898
rect 470874 401454 471194 401486
rect 470874 401218 470916 401454
rect 471152 401218 471194 401454
rect 470874 401134 471194 401218
rect 470874 400898 470916 401134
rect 471152 400898 471194 401134
rect 470874 400866 471194 400898
rect 476805 401454 477125 401486
rect 476805 401218 476847 401454
rect 477083 401218 477125 401454
rect 476805 401134 477125 401218
rect 476805 400898 476847 401134
rect 477083 400898 477125 401134
rect 476805 400866 477125 400898
rect 498874 401454 499194 401486
rect 498874 401218 498916 401454
rect 499152 401218 499194 401454
rect 498874 401134 499194 401218
rect 498874 400898 498916 401134
rect 499152 400898 499194 401134
rect 498874 400866 499194 400898
rect 504805 401454 505125 401486
rect 504805 401218 504847 401454
rect 505083 401218 505125 401454
rect 504805 401134 505125 401218
rect 504805 400898 504847 401134
rect 505083 400898 505125 401134
rect 504805 400866 505125 400898
rect 526874 401454 527194 401486
rect 526874 401218 526916 401454
rect 527152 401218 527194 401454
rect 526874 401134 527194 401218
rect 526874 400898 526916 401134
rect 527152 400898 527194 401134
rect 526874 400866 527194 400898
rect 532805 401454 533125 401486
rect 532805 401218 532847 401454
rect 533083 401218 533125 401454
rect 532805 401134 533125 401218
rect 532805 400898 532847 401134
rect 533083 400898 533125 401134
rect 532805 400866 533125 400898
rect 554874 401454 555194 401486
rect 554874 401218 554916 401454
rect 555152 401218 555194 401454
rect 554874 401134 555194 401218
rect 554874 400898 554916 401134
rect 555152 400898 555194 401134
rect 554874 400866 555194 400898
rect 560805 401454 561125 401486
rect 560805 401218 560847 401454
rect 561083 401218 561125 401454
rect 560805 401134 561125 401218
rect 560805 400898 560847 401134
rect 561083 400898 561125 401134
rect 560805 400866 561125 400898
rect -2006 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 -1386 377829
rect -2006 377509 -1386 377593
rect -2006 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 -1386 377509
rect -2006 350829 -1386 377273
rect 19910 377829 20230 377861
rect 19910 377593 19952 377829
rect 20188 377593 20230 377829
rect 19910 377509 20230 377593
rect 19910 377273 19952 377509
rect 20188 377273 20230 377509
rect 19910 377241 20230 377273
rect 25840 377829 26160 377861
rect 25840 377593 25882 377829
rect 26118 377593 26160 377829
rect 25840 377509 26160 377593
rect 25840 377273 25882 377509
rect 26118 377273 26160 377509
rect 25840 377241 26160 377273
rect 31771 377829 32091 377861
rect 31771 377593 31813 377829
rect 32049 377593 32091 377829
rect 31771 377509 32091 377593
rect 31771 377273 31813 377509
rect 32049 377273 32091 377509
rect 31771 377241 32091 377273
rect 47910 377829 48230 377861
rect 47910 377593 47952 377829
rect 48188 377593 48230 377829
rect 47910 377509 48230 377593
rect 47910 377273 47952 377509
rect 48188 377273 48230 377509
rect 47910 377241 48230 377273
rect 53840 377829 54160 377861
rect 53840 377593 53882 377829
rect 54118 377593 54160 377829
rect 53840 377509 54160 377593
rect 53840 377273 53882 377509
rect 54118 377273 54160 377509
rect 53840 377241 54160 377273
rect 59771 377829 60091 377861
rect 59771 377593 59813 377829
rect 60049 377593 60091 377829
rect 59771 377509 60091 377593
rect 59771 377273 59813 377509
rect 60049 377273 60091 377509
rect 59771 377241 60091 377273
rect 75910 377829 76230 377861
rect 75910 377593 75952 377829
rect 76188 377593 76230 377829
rect 75910 377509 76230 377593
rect 75910 377273 75952 377509
rect 76188 377273 76230 377509
rect 75910 377241 76230 377273
rect 81840 377829 82160 377861
rect 81840 377593 81882 377829
rect 82118 377593 82160 377829
rect 81840 377509 82160 377593
rect 81840 377273 81882 377509
rect 82118 377273 82160 377509
rect 81840 377241 82160 377273
rect 87771 377829 88091 377861
rect 87771 377593 87813 377829
rect 88049 377593 88091 377829
rect 87771 377509 88091 377593
rect 87771 377273 87813 377509
rect 88049 377273 88091 377509
rect 87771 377241 88091 377273
rect 103910 377829 104230 377861
rect 103910 377593 103952 377829
rect 104188 377593 104230 377829
rect 103910 377509 104230 377593
rect 103910 377273 103952 377509
rect 104188 377273 104230 377509
rect 103910 377241 104230 377273
rect 109840 377829 110160 377861
rect 109840 377593 109882 377829
rect 110118 377593 110160 377829
rect 109840 377509 110160 377593
rect 109840 377273 109882 377509
rect 110118 377273 110160 377509
rect 109840 377241 110160 377273
rect 115771 377829 116091 377861
rect 115771 377593 115813 377829
rect 116049 377593 116091 377829
rect 115771 377509 116091 377593
rect 115771 377273 115813 377509
rect 116049 377273 116091 377509
rect 115771 377241 116091 377273
rect 131910 377829 132230 377861
rect 131910 377593 131952 377829
rect 132188 377593 132230 377829
rect 131910 377509 132230 377593
rect 131910 377273 131952 377509
rect 132188 377273 132230 377509
rect 131910 377241 132230 377273
rect 137840 377829 138160 377861
rect 137840 377593 137882 377829
rect 138118 377593 138160 377829
rect 137840 377509 138160 377593
rect 137840 377273 137882 377509
rect 138118 377273 138160 377509
rect 137840 377241 138160 377273
rect 143771 377829 144091 377861
rect 143771 377593 143813 377829
rect 144049 377593 144091 377829
rect 143771 377509 144091 377593
rect 143771 377273 143813 377509
rect 144049 377273 144091 377509
rect 143771 377241 144091 377273
rect 159910 377829 160230 377861
rect 159910 377593 159952 377829
rect 160188 377593 160230 377829
rect 159910 377509 160230 377593
rect 159910 377273 159952 377509
rect 160188 377273 160230 377509
rect 159910 377241 160230 377273
rect 165840 377829 166160 377861
rect 165840 377593 165882 377829
rect 166118 377593 166160 377829
rect 165840 377509 166160 377593
rect 165840 377273 165882 377509
rect 166118 377273 166160 377509
rect 165840 377241 166160 377273
rect 171771 377829 172091 377861
rect 171771 377593 171813 377829
rect 172049 377593 172091 377829
rect 171771 377509 172091 377593
rect 171771 377273 171813 377509
rect 172049 377273 172091 377509
rect 171771 377241 172091 377273
rect 187910 377829 188230 377861
rect 187910 377593 187952 377829
rect 188188 377593 188230 377829
rect 187910 377509 188230 377593
rect 187910 377273 187952 377509
rect 188188 377273 188230 377509
rect 187910 377241 188230 377273
rect 193840 377829 194160 377861
rect 193840 377593 193882 377829
rect 194118 377593 194160 377829
rect 193840 377509 194160 377593
rect 193840 377273 193882 377509
rect 194118 377273 194160 377509
rect 193840 377241 194160 377273
rect 199771 377829 200091 377861
rect 199771 377593 199813 377829
rect 200049 377593 200091 377829
rect 199771 377509 200091 377593
rect 199771 377273 199813 377509
rect 200049 377273 200091 377509
rect 199771 377241 200091 377273
rect 215910 377829 216230 377861
rect 215910 377593 215952 377829
rect 216188 377593 216230 377829
rect 215910 377509 216230 377593
rect 215910 377273 215952 377509
rect 216188 377273 216230 377509
rect 215910 377241 216230 377273
rect 221840 377829 222160 377861
rect 221840 377593 221882 377829
rect 222118 377593 222160 377829
rect 221840 377509 222160 377593
rect 221840 377273 221882 377509
rect 222118 377273 222160 377509
rect 221840 377241 222160 377273
rect 227771 377829 228091 377861
rect 227771 377593 227813 377829
rect 228049 377593 228091 377829
rect 227771 377509 228091 377593
rect 227771 377273 227813 377509
rect 228049 377273 228091 377509
rect 227771 377241 228091 377273
rect 243910 377829 244230 377861
rect 243910 377593 243952 377829
rect 244188 377593 244230 377829
rect 243910 377509 244230 377593
rect 243910 377273 243952 377509
rect 244188 377273 244230 377509
rect 243910 377241 244230 377273
rect 249840 377829 250160 377861
rect 249840 377593 249882 377829
rect 250118 377593 250160 377829
rect 249840 377509 250160 377593
rect 249840 377273 249882 377509
rect 250118 377273 250160 377509
rect 249840 377241 250160 377273
rect 255771 377829 256091 377861
rect 255771 377593 255813 377829
rect 256049 377593 256091 377829
rect 255771 377509 256091 377593
rect 255771 377273 255813 377509
rect 256049 377273 256091 377509
rect 255771 377241 256091 377273
rect 271910 377829 272230 377861
rect 271910 377593 271952 377829
rect 272188 377593 272230 377829
rect 271910 377509 272230 377593
rect 271910 377273 271952 377509
rect 272188 377273 272230 377509
rect 271910 377241 272230 377273
rect 277840 377829 278160 377861
rect 277840 377593 277882 377829
rect 278118 377593 278160 377829
rect 277840 377509 278160 377593
rect 277840 377273 277882 377509
rect 278118 377273 278160 377509
rect 277840 377241 278160 377273
rect 283771 377829 284091 377861
rect 283771 377593 283813 377829
rect 284049 377593 284091 377829
rect 283771 377509 284091 377593
rect 283771 377273 283813 377509
rect 284049 377273 284091 377509
rect 283771 377241 284091 377273
rect 299910 377829 300230 377861
rect 299910 377593 299952 377829
rect 300188 377593 300230 377829
rect 299910 377509 300230 377593
rect 299910 377273 299952 377509
rect 300188 377273 300230 377509
rect 299910 377241 300230 377273
rect 305840 377829 306160 377861
rect 305840 377593 305882 377829
rect 306118 377593 306160 377829
rect 305840 377509 306160 377593
rect 305840 377273 305882 377509
rect 306118 377273 306160 377509
rect 305840 377241 306160 377273
rect 311771 377829 312091 377861
rect 311771 377593 311813 377829
rect 312049 377593 312091 377829
rect 311771 377509 312091 377593
rect 311771 377273 311813 377509
rect 312049 377273 312091 377509
rect 311771 377241 312091 377273
rect 327910 377829 328230 377861
rect 327910 377593 327952 377829
rect 328188 377593 328230 377829
rect 327910 377509 328230 377593
rect 327910 377273 327952 377509
rect 328188 377273 328230 377509
rect 327910 377241 328230 377273
rect 333840 377829 334160 377861
rect 333840 377593 333882 377829
rect 334118 377593 334160 377829
rect 333840 377509 334160 377593
rect 333840 377273 333882 377509
rect 334118 377273 334160 377509
rect 333840 377241 334160 377273
rect 339771 377829 340091 377861
rect 339771 377593 339813 377829
rect 340049 377593 340091 377829
rect 339771 377509 340091 377593
rect 339771 377273 339813 377509
rect 340049 377273 340091 377509
rect 339771 377241 340091 377273
rect 355910 377829 356230 377861
rect 355910 377593 355952 377829
rect 356188 377593 356230 377829
rect 355910 377509 356230 377593
rect 355910 377273 355952 377509
rect 356188 377273 356230 377509
rect 355910 377241 356230 377273
rect 361840 377829 362160 377861
rect 361840 377593 361882 377829
rect 362118 377593 362160 377829
rect 361840 377509 362160 377593
rect 361840 377273 361882 377509
rect 362118 377273 362160 377509
rect 361840 377241 362160 377273
rect 367771 377829 368091 377861
rect 367771 377593 367813 377829
rect 368049 377593 368091 377829
rect 367771 377509 368091 377593
rect 367771 377273 367813 377509
rect 368049 377273 368091 377509
rect 367771 377241 368091 377273
rect 383910 377829 384230 377861
rect 383910 377593 383952 377829
rect 384188 377593 384230 377829
rect 383910 377509 384230 377593
rect 383910 377273 383952 377509
rect 384188 377273 384230 377509
rect 383910 377241 384230 377273
rect 389840 377829 390160 377861
rect 389840 377593 389882 377829
rect 390118 377593 390160 377829
rect 389840 377509 390160 377593
rect 389840 377273 389882 377509
rect 390118 377273 390160 377509
rect 389840 377241 390160 377273
rect 395771 377829 396091 377861
rect 395771 377593 395813 377829
rect 396049 377593 396091 377829
rect 395771 377509 396091 377593
rect 395771 377273 395813 377509
rect 396049 377273 396091 377509
rect 395771 377241 396091 377273
rect 411910 377829 412230 377861
rect 411910 377593 411952 377829
rect 412188 377593 412230 377829
rect 411910 377509 412230 377593
rect 411910 377273 411952 377509
rect 412188 377273 412230 377509
rect 411910 377241 412230 377273
rect 417840 377829 418160 377861
rect 417840 377593 417882 377829
rect 418118 377593 418160 377829
rect 417840 377509 418160 377593
rect 417840 377273 417882 377509
rect 418118 377273 418160 377509
rect 417840 377241 418160 377273
rect 423771 377829 424091 377861
rect 423771 377593 423813 377829
rect 424049 377593 424091 377829
rect 423771 377509 424091 377593
rect 423771 377273 423813 377509
rect 424049 377273 424091 377509
rect 423771 377241 424091 377273
rect 439910 377829 440230 377861
rect 439910 377593 439952 377829
rect 440188 377593 440230 377829
rect 439910 377509 440230 377593
rect 439910 377273 439952 377509
rect 440188 377273 440230 377509
rect 439910 377241 440230 377273
rect 445840 377829 446160 377861
rect 445840 377593 445882 377829
rect 446118 377593 446160 377829
rect 445840 377509 446160 377593
rect 445840 377273 445882 377509
rect 446118 377273 446160 377509
rect 445840 377241 446160 377273
rect 451771 377829 452091 377861
rect 451771 377593 451813 377829
rect 452049 377593 452091 377829
rect 451771 377509 452091 377593
rect 451771 377273 451813 377509
rect 452049 377273 452091 377509
rect 451771 377241 452091 377273
rect 467910 377829 468230 377861
rect 467910 377593 467952 377829
rect 468188 377593 468230 377829
rect 467910 377509 468230 377593
rect 467910 377273 467952 377509
rect 468188 377273 468230 377509
rect 467910 377241 468230 377273
rect 473840 377829 474160 377861
rect 473840 377593 473882 377829
rect 474118 377593 474160 377829
rect 473840 377509 474160 377593
rect 473840 377273 473882 377509
rect 474118 377273 474160 377509
rect 473840 377241 474160 377273
rect 479771 377829 480091 377861
rect 479771 377593 479813 377829
rect 480049 377593 480091 377829
rect 479771 377509 480091 377593
rect 479771 377273 479813 377509
rect 480049 377273 480091 377509
rect 479771 377241 480091 377273
rect 495910 377829 496230 377861
rect 495910 377593 495952 377829
rect 496188 377593 496230 377829
rect 495910 377509 496230 377593
rect 495910 377273 495952 377509
rect 496188 377273 496230 377509
rect 495910 377241 496230 377273
rect 501840 377829 502160 377861
rect 501840 377593 501882 377829
rect 502118 377593 502160 377829
rect 501840 377509 502160 377593
rect 501840 377273 501882 377509
rect 502118 377273 502160 377509
rect 501840 377241 502160 377273
rect 507771 377829 508091 377861
rect 507771 377593 507813 377829
rect 508049 377593 508091 377829
rect 507771 377509 508091 377593
rect 507771 377273 507813 377509
rect 508049 377273 508091 377509
rect 507771 377241 508091 377273
rect 523910 377829 524230 377861
rect 523910 377593 523952 377829
rect 524188 377593 524230 377829
rect 523910 377509 524230 377593
rect 523910 377273 523952 377509
rect 524188 377273 524230 377509
rect 523910 377241 524230 377273
rect 529840 377829 530160 377861
rect 529840 377593 529882 377829
rect 530118 377593 530160 377829
rect 529840 377509 530160 377593
rect 529840 377273 529882 377509
rect 530118 377273 530160 377509
rect 529840 377241 530160 377273
rect 535771 377829 536091 377861
rect 535771 377593 535813 377829
rect 536049 377593 536091 377829
rect 535771 377509 536091 377593
rect 535771 377273 535813 377509
rect 536049 377273 536091 377509
rect 535771 377241 536091 377273
rect 551910 377829 552230 377861
rect 551910 377593 551952 377829
rect 552188 377593 552230 377829
rect 551910 377509 552230 377593
rect 551910 377273 551952 377509
rect 552188 377273 552230 377509
rect 551910 377241 552230 377273
rect 557840 377829 558160 377861
rect 557840 377593 557882 377829
rect 558118 377593 558160 377829
rect 557840 377509 558160 377593
rect 557840 377273 557882 377509
rect 558118 377273 558160 377509
rect 557840 377241 558160 377273
rect 563771 377829 564091 377861
rect 563771 377593 563813 377829
rect 564049 377593 564091 377829
rect 563771 377509 564091 377593
rect 563771 377273 563813 377509
rect 564049 377273 564091 377509
rect 563771 377241 564091 377273
rect 573494 377829 574114 404273
rect 573494 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 574114 377829
rect 573494 377509 574114 377593
rect 573494 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 574114 377509
rect 22874 374454 23194 374486
rect 22874 374218 22916 374454
rect 23152 374218 23194 374454
rect 22874 374134 23194 374218
rect 22874 373898 22916 374134
rect 23152 373898 23194 374134
rect 22874 373866 23194 373898
rect 28805 374454 29125 374486
rect 28805 374218 28847 374454
rect 29083 374218 29125 374454
rect 28805 374134 29125 374218
rect 28805 373898 28847 374134
rect 29083 373898 29125 374134
rect 28805 373866 29125 373898
rect 50874 374454 51194 374486
rect 50874 374218 50916 374454
rect 51152 374218 51194 374454
rect 50874 374134 51194 374218
rect 50874 373898 50916 374134
rect 51152 373898 51194 374134
rect 50874 373866 51194 373898
rect 56805 374454 57125 374486
rect 56805 374218 56847 374454
rect 57083 374218 57125 374454
rect 56805 374134 57125 374218
rect 56805 373898 56847 374134
rect 57083 373898 57125 374134
rect 56805 373866 57125 373898
rect 78874 374454 79194 374486
rect 78874 374218 78916 374454
rect 79152 374218 79194 374454
rect 78874 374134 79194 374218
rect 78874 373898 78916 374134
rect 79152 373898 79194 374134
rect 78874 373866 79194 373898
rect 84805 374454 85125 374486
rect 84805 374218 84847 374454
rect 85083 374218 85125 374454
rect 84805 374134 85125 374218
rect 84805 373898 84847 374134
rect 85083 373898 85125 374134
rect 84805 373866 85125 373898
rect 106874 374454 107194 374486
rect 106874 374218 106916 374454
rect 107152 374218 107194 374454
rect 106874 374134 107194 374218
rect 106874 373898 106916 374134
rect 107152 373898 107194 374134
rect 106874 373866 107194 373898
rect 112805 374454 113125 374486
rect 112805 374218 112847 374454
rect 113083 374218 113125 374454
rect 112805 374134 113125 374218
rect 112805 373898 112847 374134
rect 113083 373898 113125 374134
rect 112805 373866 113125 373898
rect 134874 374454 135194 374486
rect 134874 374218 134916 374454
rect 135152 374218 135194 374454
rect 134874 374134 135194 374218
rect 134874 373898 134916 374134
rect 135152 373898 135194 374134
rect 134874 373866 135194 373898
rect 140805 374454 141125 374486
rect 140805 374218 140847 374454
rect 141083 374218 141125 374454
rect 140805 374134 141125 374218
rect 140805 373898 140847 374134
rect 141083 373898 141125 374134
rect 140805 373866 141125 373898
rect 162874 374454 163194 374486
rect 162874 374218 162916 374454
rect 163152 374218 163194 374454
rect 162874 374134 163194 374218
rect 162874 373898 162916 374134
rect 163152 373898 163194 374134
rect 162874 373866 163194 373898
rect 168805 374454 169125 374486
rect 168805 374218 168847 374454
rect 169083 374218 169125 374454
rect 168805 374134 169125 374218
rect 168805 373898 168847 374134
rect 169083 373898 169125 374134
rect 168805 373866 169125 373898
rect 190874 374454 191194 374486
rect 190874 374218 190916 374454
rect 191152 374218 191194 374454
rect 190874 374134 191194 374218
rect 190874 373898 190916 374134
rect 191152 373898 191194 374134
rect 190874 373866 191194 373898
rect 196805 374454 197125 374486
rect 196805 374218 196847 374454
rect 197083 374218 197125 374454
rect 196805 374134 197125 374218
rect 196805 373898 196847 374134
rect 197083 373898 197125 374134
rect 196805 373866 197125 373898
rect 218874 374454 219194 374486
rect 218874 374218 218916 374454
rect 219152 374218 219194 374454
rect 218874 374134 219194 374218
rect 218874 373898 218916 374134
rect 219152 373898 219194 374134
rect 218874 373866 219194 373898
rect 224805 374454 225125 374486
rect 224805 374218 224847 374454
rect 225083 374218 225125 374454
rect 224805 374134 225125 374218
rect 224805 373898 224847 374134
rect 225083 373898 225125 374134
rect 224805 373866 225125 373898
rect 246874 374454 247194 374486
rect 246874 374218 246916 374454
rect 247152 374218 247194 374454
rect 246874 374134 247194 374218
rect 246874 373898 246916 374134
rect 247152 373898 247194 374134
rect 246874 373866 247194 373898
rect 252805 374454 253125 374486
rect 252805 374218 252847 374454
rect 253083 374218 253125 374454
rect 252805 374134 253125 374218
rect 252805 373898 252847 374134
rect 253083 373898 253125 374134
rect 252805 373866 253125 373898
rect 274874 374454 275194 374486
rect 274874 374218 274916 374454
rect 275152 374218 275194 374454
rect 274874 374134 275194 374218
rect 274874 373898 274916 374134
rect 275152 373898 275194 374134
rect 274874 373866 275194 373898
rect 280805 374454 281125 374486
rect 280805 374218 280847 374454
rect 281083 374218 281125 374454
rect 280805 374134 281125 374218
rect 280805 373898 280847 374134
rect 281083 373898 281125 374134
rect 280805 373866 281125 373898
rect 302874 374454 303194 374486
rect 302874 374218 302916 374454
rect 303152 374218 303194 374454
rect 302874 374134 303194 374218
rect 302874 373898 302916 374134
rect 303152 373898 303194 374134
rect 302874 373866 303194 373898
rect 308805 374454 309125 374486
rect 308805 374218 308847 374454
rect 309083 374218 309125 374454
rect 308805 374134 309125 374218
rect 308805 373898 308847 374134
rect 309083 373898 309125 374134
rect 308805 373866 309125 373898
rect 330874 374454 331194 374486
rect 330874 374218 330916 374454
rect 331152 374218 331194 374454
rect 330874 374134 331194 374218
rect 330874 373898 330916 374134
rect 331152 373898 331194 374134
rect 330874 373866 331194 373898
rect 336805 374454 337125 374486
rect 336805 374218 336847 374454
rect 337083 374218 337125 374454
rect 336805 374134 337125 374218
rect 336805 373898 336847 374134
rect 337083 373898 337125 374134
rect 336805 373866 337125 373898
rect 358874 374454 359194 374486
rect 358874 374218 358916 374454
rect 359152 374218 359194 374454
rect 358874 374134 359194 374218
rect 358874 373898 358916 374134
rect 359152 373898 359194 374134
rect 358874 373866 359194 373898
rect 364805 374454 365125 374486
rect 364805 374218 364847 374454
rect 365083 374218 365125 374454
rect 364805 374134 365125 374218
rect 364805 373898 364847 374134
rect 365083 373898 365125 374134
rect 364805 373866 365125 373898
rect 386874 374454 387194 374486
rect 386874 374218 386916 374454
rect 387152 374218 387194 374454
rect 386874 374134 387194 374218
rect 386874 373898 386916 374134
rect 387152 373898 387194 374134
rect 386874 373866 387194 373898
rect 392805 374454 393125 374486
rect 392805 374218 392847 374454
rect 393083 374218 393125 374454
rect 392805 374134 393125 374218
rect 392805 373898 392847 374134
rect 393083 373898 393125 374134
rect 392805 373866 393125 373898
rect 414874 374454 415194 374486
rect 414874 374218 414916 374454
rect 415152 374218 415194 374454
rect 414874 374134 415194 374218
rect 414874 373898 414916 374134
rect 415152 373898 415194 374134
rect 414874 373866 415194 373898
rect 420805 374454 421125 374486
rect 420805 374218 420847 374454
rect 421083 374218 421125 374454
rect 420805 374134 421125 374218
rect 420805 373898 420847 374134
rect 421083 373898 421125 374134
rect 420805 373866 421125 373898
rect 442874 374454 443194 374486
rect 442874 374218 442916 374454
rect 443152 374218 443194 374454
rect 442874 374134 443194 374218
rect 442874 373898 442916 374134
rect 443152 373898 443194 374134
rect 442874 373866 443194 373898
rect 448805 374454 449125 374486
rect 448805 374218 448847 374454
rect 449083 374218 449125 374454
rect 448805 374134 449125 374218
rect 448805 373898 448847 374134
rect 449083 373898 449125 374134
rect 448805 373866 449125 373898
rect 470874 374454 471194 374486
rect 470874 374218 470916 374454
rect 471152 374218 471194 374454
rect 470874 374134 471194 374218
rect 470874 373898 470916 374134
rect 471152 373898 471194 374134
rect 470874 373866 471194 373898
rect 476805 374454 477125 374486
rect 476805 374218 476847 374454
rect 477083 374218 477125 374454
rect 476805 374134 477125 374218
rect 476805 373898 476847 374134
rect 477083 373898 477125 374134
rect 476805 373866 477125 373898
rect 498874 374454 499194 374486
rect 498874 374218 498916 374454
rect 499152 374218 499194 374454
rect 498874 374134 499194 374218
rect 498874 373898 498916 374134
rect 499152 373898 499194 374134
rect 498874 373866 499194 373898
rect 504805 374454 505125 374486
rect 504805 374218 504847 374454
rect 505083 374218 505125 374454
rect 504805 374134 505125 374218
rect 504805 373898 504847 374134
rect 505083 373898 505125 374134
rect 504805 373866 505125 373898
rect 526874 374454 527194 374486
rect 526874 374218 526916 374454
rect 527152 374218 527194 374454
rect 526874 374134 527194 374218
rect 526874 373898 526916 374134
rect 527152 373898 527194 374134
rect 526874 373866 527194 373898
rect 532805 374454 533125 374486
rect 532805 374218 532847 374454
rect 533083 374218 533125 374454
rect 532805 374134 533125 374218
rect 532805 373898 532847 374134
rect 533083 373898 533125 374134
rect 532805 373866 533125 373898
rect 554874 374454 555194 374486
rect 554874 374218 554916 374454
rect 555152 374218 555194 374454
rect 554874 374134 555194 374218
rect 554874 373898 554916 374134
rect 555152 373898 555194 374134
rect 554874 373866 555194 373898
rect 560805 374454 561125 374486
rect 560805 374218 560847 374454
rect 561083 374218 561125 374454
rect 560805 374134 561125 374218
rect 560805 373898 560847 374134
rect 561083 373898 561125 374134
rect 560805 373866 561125 373898
rect -2006 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 -1386 350829
rect -2006 350509 -1386 350593
rect -2006 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 -1386 350509
rect -2006 323829 -1386 350273
rect 19910 350829 20230 350861
rect 19910 350593 19952 350829
rect 20188 350593 20230 350829
rect 19910 350509 20230 350593
rect 19910 350273 19952 350509
rect 20188 350273 20230 350509
rect 19910 350241 20230 350273
rect 25840 350829 26160 350861
rect 25840 350593 25882 350829
rect 26118 350593 26160 350829
rect 25840 350509 26160 350593
rect 25840 350273 25882 350509
rect 26118 350273 26160 350509
rect 25840 350241 26160 350273
rect 31771 350829 32091 350861
rect 31771 350593 31813 350829
rect 32049 350593 32091 350829
rect 31771 350509 32091 350593
rect 31771 350273 31813 350509
rect 32049 350273 32091 350509
rect 31771 350241 32091 350273
rect 47910 350829 48230 350861
rect 47910 350593 47952 350829
rect 48188 350593 48230 350829
rect 47910 350509 48230 350593
rect 47910 350273 47952 350509
rect 48188 350273 48230 350509
rect 47910 350241 48230 350273
rect 53840 350829 54160 350861
rect 53840 350593 53882 350829
rect 54118 350593 54160 350829
rect 53840 350509 54160 350593
rect 53840 350273 53882 350509
rect 54118 350273 54160 350509
rect 53840 350241 54160 350273
rect 59771 350829 60091 350861
rect 59771 350593 59813 350829
rect 60049 350593 60091 350829
rect 59771 350509 60091 350593
rect 59771 350273 59813 350509
rect 60049 350273 60091 350509
rect 59771 350241 60091 350273
rect 75910 350829 76230 350861
rect 75910 350593 75952 350829
rect 76188 350593 76230 350829
rect 75910 350509 76230 350593
rect 75910 350273 75952 350509
rect 76188 350273 76230 350509
rect 75910 350241 76230 350273
rect 81840 350829 82160 350861
rect 81840 350593 81882 350829
rect 82118 350593 82160 350829
rect 81840 350509 82160 350593
rect 81840 350273 81882 350509
rect 82118 350273 82160 350509
rect 81840 350241 82160 350273
rect 87771 350829 88091 350861
rect 87771 350593 87813 350829
rect 88049 350593 88091 350829
rect 87771 350509 88091 350593
rect 87771 350273 87813 350509
rect 88049 350273 88091 350509
rect 87771 350241 88091 350273
rect 103910 350829 104230 350861
rect 103910 350593 103952 350829
rect 104188 350593 104230 350829
rect 103910 350509 104230 350593
rect 103910 350273 103952 350509
rect 104188 350273 104230 350509
rect 103910 350241 104230 350273
rect 109840 350829 110160 350861
rect 109840 350593 109882 350829
rect 110118 350593 110160 350829
rect 109840 350509 110160 350593
rect 109840 350273 109882 350509
rect 110118 350273 110160 350509
rect 109840 350241 110160 350273
rect 115771 350829 116091 350861
rect 115771 350593 115813 350829
rect 116049 350593 116091 350829
rect 115771 350509 116091 350593
rect 115771 350273 115813 350509
rect 116049 350273 116091 350509
rect 115771 350241 116091 350273
rect 131910 350829 132230 350861
rect 131910 350593 131952 350829
rect 132188 350593 132230 350829
rect 131910 350509 132230 350593
rect 131910 350273 131952 350509
rect 132188 350273 132230 350509
rect 131910 350241 132230 350273
rect 137840 350829 138160 350861
rect 137840 350593 137882 350829
rect 138118 350593 138160 350829
rect 137840 350509 138160 350593
rect 137840 350273 137882 350509
rect 138118 350273 138160 350509
rect 137840 350241 138160 350273
rect 143771 350829 144091 350861
rect 143771 350593 143813 350829
rect 144049 350593 144091 350829
rect 143771 350509 144091 350593
rect 143771 350273 143813 350509
rect 144049 350273 144091 350509
rect 143771 350241 144091 350273
rect 159910 350829 160230 350861
rect 159910 350593 159952 350829
rect 160188 350593 160230 350829
rect 159910 350509 160230 350593
rect 159910 350273 159952 350509
rect 160188 350273 160230 350509
rect 159910 350241 160230 350273
rect 165840 350829 166160 350861
rect 165840 350593 165882 350829
rect 166118 350593 166160 350829
rect 165840 350509 166160 350593
rect 165840 350273 165882 350509
rect 166118 350273 166160 350509
rect 165840 350241 166160 350273
rect 171771 350829 172091 350861
rect 171771 350593 171813 350829
rect 172049 350593 172091 350829
rect 171771 350509 172091 350593
rect 171771 350273 171813 350509
rect 172049 350273 172091 350509
rect 171771 350241 172091 350273
rect 187910 350829 188230 350861
rect 187910 350593 187952 350829
rect 188188 350593 188230 350829
rect 187910 350509 188230 350593
rect 187910 350273 187952 350509
rect 188188 350273 188230 350509
rect 187910 350241 188230 350273
rect 193840 350829 194160 350861
rect 193840 350593 193882 350829
rect 194118 350593 194160 350829
rect 193840 350509 194160 350593
rect 193840 350273 193882 350509
rect 194118 350273 194160 350509
rect 193840 350241 194160 350273
rect 199771 350829 200091 350861
rect 199771 350593 199813 350829
rect 200049 350593 200091 350829
rect 199771 350509 200091 350593
rect 199771 350273 199813 350509
rect 200049 350273 200091 350509
rect 199771 350241 200091 350273
rect 215910 350829 216230 350861
rect 215910 350593 215952 350829
rect 216188 350593 216230 350829
rect 215910 350509 216230 350593
rect 215910 350273 215952 350509
rect 216188 350273 216230 350509
rect 215910 350241 216230 350273
rect 221840 350829 222160 350861
rect 221840 350593 221882 350829
rect 222118 350593 222160 350829
rect 221840 350509 222160 350593
rect 221840 350273 221882 350509
rect 222118 350273 222160 350509
rect 221840 350241 222160 350273
rect 227771 350829 228091 350861
rect 227771 350593 227813 350829
rect 228049 350593 228091 350829
rect 227771 350509 228091 350593
rect 227771 350273 227813 350509
rect 228049 350273 228091 350509
rect 227771 350241 228091 350273
rect 243910 350829 244230 350861
rect 243910 350593 243952 350829
rect 244188 350593 244230 350829
rect 243910 350509 244230 350593
rect 243910 350273 243952 350509
rect 244188 350273 244230 350509
rect 243910 350241 244230 350273
rect 249840 350829 250160 350861
rect 249840 350593 249882 350829
rect 250118 350593 250160 350829
rect 249840 350509 250160 350593
rect 249840 350273 249882 350509
rect 250118 350273 250160 350509
rect 249840 350241 250160 350273
rect 255771 350829 256091 350861
rect 255771 350593 255813 350829
rect 256049 350593 256091 350829
rect 255771 350509 256091 350593
rect 255771 350273 255813 350509
rect 256049 350273 256091 350509
rect 255771 350241 256091 350273
rect 271910 350829 272230 350861
rect 271910 350593 271952 350829
rect 272188 350593 272230 350829
rect 271910 350509 272230 350593
rect 271910 350273 271952 350509
rect 272188 350273 272230 350509
rect 271910 350241 272230 350273
rect 277840 350829 278160 350861
rect 277840 350593 277882 350829
rect 278118 350593 278160 350829
rect 277840 350509 278160 350593
rect 277840 350273 277882 350509
rect 278118 350273 278160 350509
rect 277840 350241 278160 350273
rect 283771 350829 284091 350861
rect 283771 350593 283813 350829
rect 284049 350593 284091 350829
rect 283771 350509 284091 350593
rect 283771 350273 283813 350509
rect 284049 350273 284091 350509
rect 283771 350241 284091 350273
rect 299910 350829 300230 350861
rect 299910 350593 299952 350829
rect 300188 350593 300230 350829
rect 299910 350509 300230 350593
rect 299910 350273 299952 350509
rect 300188 350273 300230 350509
rect 299910 350241 300230 350273
rect 305840 350829 306160 350861
rect 305840 350593 305882 350829
rect 306118 350593 306160 350829
rect 305840 350509 306160 350593
rect 305840 350273 305882 350509
rect 306118 350273 306160 350509
rect 305840 350241 306160 350273
rect 311771 350829 312091 350861
rect 311771 350593 311813 350829
rect 312049 350593 312091 350829
rect 311771 350509 312091 350593
rect 311771 350273 311813 350509
rect 312049 350273 312091 350509
rect 311771 350241 312091 350273
rect 327910 350829 328230 350861
rect 327910 350593 327952 350829
rect 328188 350593 328230 350829
rect 327910 350509 328230 350593
rect 327910 350273 327952 350509
rect 328188 350273 328230 350509
rect 327910 350241 328230 350273
rect 333840 350829 334160 350861
rect 333840 350593 333882 350829
rect 334118 350593 334160 350829
rect 333840 350509 334160 350593
rect 333840 350273 333882 350509
rect 334118 350273 334160 350509
rect 333840 350241 334160 350273
rect 339771 350829 340091 350861
rect 339771 350593 339813 350829
rect 340049 350593 340091 350829
rect 339771 350509 340091 350593
rect 339771 350273 339813 350509
rect 340049 350273 340091 350509
rect 339771 350241 340091 350273
rect 355910 350829 356230 350861
rect 355910 350593 355952 350829
rect 356188 350593 356230 350829
rect 355910 350509 356230 350593
rect 355910 350273 355952 350509
rect 356188 350273 356230 350509
rect 355910 350241 356230 350273
rect 361840 350829 362160 350861
rect 361840 350593 361882 350829
rect 362118 350593 362160 350829
rect 361840 350509 362160 350593
rect 361840 350273 361882 350509
rect 362118 350273 362160 350509
rect 361840 350241 362160 350273
rect 367771 350829 368091 350861
rect 367771 350593 367813 350829
rect 368049 350593 368091 350829
rect 367771 350509 368091 350593
rect 367771 350273 367813 350509
rect 368049 350273 368091 350509
rect 367771 350241 368091 350273
rect 383910 350829 384230 350861
rect 383910 350593 383952 350829
rect 384188 350593 384230 350829
rect 383910 350509 384230 350593
rect 383910 350273 383952 350509
rect 384188 350273 384230 350509
rect 383910 350241 384230 350273
rect 389840 350829 390160 350861
rect 389840 350593 389882 350829
rect 390118 350593 390160 350829
rect 389840 350509 390160 350593
rect 389840 350273 389882 350509
rect 390118 350273 390160 350509
rect 389840 350241 390160 350273
rect 395771 350829 396091 350861
rect 395771 350593 395813 350829
rect 396049 350593 396091 350829
rect 395771 350509 396091 350593
rect 395771 350273 395813 350509
rect 396049 350273 396091 350509
rect 395771 350241 396091 350273
rect 411910 350829 412230 350861
rect 411910 350593 411952 350829
rect 412188 350593 412230 350829
rect 411910 350509 412230 350593
rect 411910 350273 411952 350509
rect 412188 350273 412230 350509
rect 411910 350241 412230 350273
rect 417840 350829 418160 350861
rect 417840 350593 417882 350829
rect 418118 350593 418160 350829
rect 417840 350509 418160 350593
rect 417840 350273 417882 350509
rect 418118 350273 418160 350509
rect 417840 350241 418160 350273
rect 423771 350829 424091 350861
rect 423771 350593 423813 350829
rect 424049 350593 424091 350829
rect 423771 350509 424091 350593
rect 423771 350273 423813 350509
rect 424049 350273 424091 350509
rect 423771 350241 424091 350273
rect 439910 350829 440230 350861
rect 439910 350593 439952 350829
rect 440188 350593 440230 350829
rect 439910 350509 440230 350593
rect 439910 350273 439952 350509
rect 440188 350273 440230 350509
rect 439910 350241 440230 350273
rect 445840 350829 446160 350861
rect 445840 350593 445882 350829
rect 446118 350593 446160 350829
rect 445840 350509 446160 350593
rect 445840 350273 445882 350509
rect 446118 350273 446160 350509
rect 445840 350241 446160 350273
rect 451771 350829 452091 350861
rect 451771 350593 451813 350829
rect 452049 350593 452091 350829
rect 451771 350509 452091 350593
rect 451771 350273 451813 350509
rect 452049 350273 452091 350509
rect 451771 350241 452091 350273
rect 467910 350829 468230 350861
rect 467910 350593 467952 350829
rect 468188 350593 468230 350829
rect 467910 350509 468230 350593
rect 467910 350273 467952 350509
rect 468188 350273 468230 350509
rect 467910 350241 468230 350273
rect 473840 350829 474160 350861
rect 473840 350593 473882 350829
rect 474118 350593 474160 350829
rect 473840 350509 474160 350593
rect 473840 350273 473882 350509
rect 474118 350273 474160 350509
rect 473840 350241 474160 350273
rect 479771 350829 480091 350861
rect 479771 350593 479813 350829
rect 480049 350593 480091 350829
rect 479771 350509 480091 350593
rect 479771 350273 479813 350509
rect 480049 350273 480091 350509
rect 479771 350241 480091 350273
rect 495910 350829 496230 350861
rect 495910 350593 495952 350829
rect 496188 350593 496230 350829
rect 495910 350509 496230 350593
rect 495910 350273 495952 350509
rect 496188 350273 496230 350509
rect 495910 350241 496230 350273
rect 501840 350829 502160 350861
rect 501840 350593 501882 350829
rect 502118 350593 502160 350829
rect 501840 350509 502160 350593
rect 501840 350273 501882 350509
rect 502118 350273 502160 350509
rect 501840 350241 502160 350273
rect 507771 350829 508091 350861
rect 507771 350593 507813 350829
rect 508049 350593 508091 350829
rect 507771 350509 508091 350593
rect 507771 350273 507813 350509
rect 508049 350273 508091 350509
rect 507771 350241 508091 350273
rect 523910 350829 524230 350861
rect 523910 350593 523952 350829
rect 524188 350593 524230 350829
rect 523910 350509 524230 350593
rect 523910 350273 523952 350509
rect 524188 350273 524230 350509
rect 523910 350241 524230 350273
rect 529840 350829 530160 350861
rect 529840 350593 529882 350829
rect 530118 350593 530160 350829
rect 529840 350509 530160 350593
rect 529840 350273 529882 350509
rect 530118 350273 530160 350509
rect 529840 350241 530160 350273
rect 535771 350829 536091 350861
rect 535771 350593 535813 350829
rect 536049 350593 536091 350829
rect 535771 350509 536091 350593
rect 535771 350273 535813 350509
rect 536049 350273 536091 350509
rect 535771 350241 536091 350273
rect 551910 350829 552230 350861
rect 551910 350593 551952 350829
rect 552188 350593 552230 350829
rect 551910 350509 552230 350593
rect 551910 350273 551952 350509
rect 552188 350273 552230 350509
rect 551910 350241 552230 350273
rect 557840 350829 558160 350861
rect 557840 350593 557882 350829
rect 558118 350593 558160 350829
rect 557840 350509 558160 350593
rect 557840 350273 557882 350509
rect 558118 350273 558160 350509
rect 557840 350241 558160 350273
rect 563771 350829 564091 350861
rect 563771 350593 563813 350829
rect 564049 350593 564091 350829
rect 563771 350509 564091 350593
rect 563771 350273 563813 350509
rect 564049 350273 564091 350509
rect 563771 350241 564091 350273
rect 573494 350829 574114 377273
rect 573494 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 574114 350829
rect 573494 350509 574114 350593
rect 573494 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 574114 350509
rect 22874 347454 23194 347486
rect 22874 347218 22916 347454
rect 23152 347218 23194 347454
rect 22874 347134 23194 347218
rect 22874 346898 22916 347134
rect 23152 346898 23194 347134
rect 22874 346866 23194 346898
rect 28805 347454 29125 347486
rect 28805 347218 28847 347454
rect 29083 347218 29125 347454
rect 28805 347134 29125 347218
rect 28805 346898 28847 347134
rect 29083 346898 29125 347134
rect 28805 346866 29125 346898
rect 50874 347454 51194 347486
rect 50874 347218 50916 347454
rect 51152 347218 51194 347454
rect 50874 347134 51194 347218
rect 50874 346898 50916 347134
rect 51152 346898 51194 347134
rect 50874 346866 51194 346898
rect 56805 347454 57125 347486
rect 56805 347218 56847 347454
rect 57083 347218 57125 347454
rect 56805 347134 57125 347218
rect 56805 346898 56847 347134
rect 57083 346898 57125 347134
rect 56805 346866 57125 346898
rect 78874 347454 79194 347486
rect 78874 347218 78916 347454
rect 79152 347218 79194 347454
rect 78874 347134 79194 347218
rect 78874 346898 78916 347134
rect 79152 346898 79194 347134
rect 78874 346866 79194 346898
rect 84805 347454 85125 347486
rect 84805 347218 84847 347454
rect 85083 347218 85125 347454
rect 84805 347134 85125 347218
rect 84805 346898 84847 347134
rect 85083 346898 85125 347134
rect 84805 346866 85125 346898
rect 106874 347454 107194 347486
rect 106874 347218 106916 347454
rect 107152 347218 107194 347454
rect 106874 347134 107194 347218
rect 106874 346898 106916 347134
rect 107152 346898 107194 347134
rect 106874 346866 107194 346898
rect 112805 347454 113125 347486
rect 112805 347218 112847 347454
rect 113083 347218 113125 347454
rect 112805 347134 113125 347218
rect 112805 346898 112847 347134
rect 113083 346898 113125 347134
rect 112805 346866 113125 346898
rect 134874 347454 135194 347486
rect 134874 347218 134916 347454
rect 135152 347218 135194 347454
rect 134874 347134 135194 347218
rect 134874 346898 134916 347134
rect 135152 346898 135194 347134
rect 134874 346866 135194 346898
rect 140805 347454 141125 347486
rect 140805 347218 140847 347454
rect 141083 347218 141125 347454
rect 140805 347134 141125 347218
rect 140805 346898 140847 347134
rect 141083 346898 141125 347134
rect 140805 346866 141125 346898
rect 162874 347454 163194 347486
rect 162874 347218 162916 347454
rect 163152 347218 163194 347454
rect 162874 347134 163194 347218
rect 162874 346898 162916 347134
rect 163152 346898 163194 347134
rect 162874 346866 163194 346898
rect 168805 347454 169125 347486
rect 168805 347218 168847 347454
rect 169083 347218 169125 347454
rect 168805 347134 169125 347218
rect 168805 346898 168847 347134
rect 169083 346898 169125 347134
rect 168805 346866 169125 346898
rect 190874 347454 191194 347486
rect 190874 347218 190916 347454
rect 191152 347218 191194 347454
rect 190874 347134 191194 347218
rect 190874 346898 190916 347134
rect 191152 346898 191194 347134
rect 190874 346866 191194 346898
rect 196805 347454 197125 347486
rect 196805 347218 196847 347454
rect 197083 347218 197125 347454
rect 196805 347134 197125 347218
rect 196805 346898 196847 347134
rect 197083 346898 197125 347134
rect 196805 346866 197125 346898
rect 218874 347454 219194 347486
rect 218874 347218 218916 347454
rect 219152 347218 219194 347454
rect 218874 347134 219194 347218
rect 218874 346898 218916 347134
rect 219152 346898 219194 347134
rect 218874 346866 219194 346898
rect 224805 347454 225125 347486
rect 224805 347218 224847 347454
rect 225083 347218 225125 347454
rect 224805 347134 225125 347218
rect 224805 346898 224847 347134
rect 225083 346898 225125 347134
rect 224805 346866 225125 346898
rect 246874 347454 247194 347486
rect 246874 347218 246916 347454
rect 247152 347218 247194 347454
rect 246874 347134 247194 347218
rect 246874 346898 246916 347134
rect 247152 346898 247194 347134
rect 246874 346866 247194 346898
rect 252805 347454 253125 347486
rect 252805 347218 252847 347454
rect 253083 347218 253125 347454
rect 252805 347134 253125 347218
rect 252805 346898 252847 347134
rect 253083 346898 253125 347134
rect 252805 346866 253125 346898
rect 274874 347454 275194 347486
rect 274874 347218 274916 347454
rect 275152 347218 275194 347454
rect 274874 347134 275194 347218
rect 274874 346898 274916 347134
rect 275152 346898 275194 347134
rect 274874 346866 275194 346898
rect 280805 347454 281125 347486
rect 280805 347218 280847 347454
rect 281083 347218 281125 347454
rect 280805 347134 281125 347218
rect 280805 346898 280847 347134
rect 281083 346898 281125 347134
rect 280805 346866 281125 346898
rect 302874 347454 303194 347486
rect 302874 347218 302916 347454
rect 303152 347218 303194 347454
rect 302874 347134 303194 347218
rect 302874 346898 302916 347134
rect 303152 346898 303194 347134
rect 302874 346866 303194 346898
rect 308805 347454 309125 347486
rect 308805 347218 308847 347454
rect 309083 347218 309125 347454
rect 308805 347134 309125 347218
rect 308805 346898 308847 347134
rect 309083 346898 309125 347134
rect 308805 346866 309125 346898
rect 330874 347454 331194 347486
rect 330874 347218 330916 347454
rect 331152 347218 331194 347454
rect 330874 347134 331194 347218
rect 330874 346898 330916 347134
rect 331152 346898 331194 347134
rect 330874 346866 331194 346898
rect 336805 347454 337125 347486
rect 336805 347218 336847 347454
rect 337083 347218 337125 347454
rect 336805 347134 337125 347218
rect 336805 346898 336847 347134
rect 337083 346898 337125 347134
rect 336805 346866 337125 346898
rect 358874 347454 359194 347486
rect 358874 347218 358916 347454
rect 359152 347218 359194 347454
rect 358874 347134 359194 347218
rect 358874 346898 358916 347134
rect 359152 346898 359194 347134
rect 358874 346866 359194 346898
rect 364805 347454 365125 347486
rect 364805 347218 364847 347454
rect 365083 347218 365125 347454
rect 364805 347134 365125 347218
rect 364805 346898 364847 347134
rect 365083 346898 365125 347134
rect 364805 346866 365125 346898
rect 386874 347454 387194 347486
rect 386874 347218 386916 347454
rect 387152 347218 387194 347454
rect 386874 347134 387194 347218
rect 386874 346898 386916 347134
rect 387152 346898 387194 347134
rect 386874 346866 387194 346898
rect 392805 347454 393125 347486
rect 392805 347218 392847 347454
rect 393083 347218 393125 347454
rect 392805 347134 393125 347218
rect 392805 346898 392847 347134
rect 393083 346898 393125 347134
rect 392805 346866 393125 346898
rect 414874 347454 415194 347486
rect 414874 347218 414916 347454
rect 415152 347218 415194 347454
rect 414874 347134 415194 347218
rect 414874 346898 414916 347134
rect 415152 346898 415194 347134
rect 414874 346866 415194 346898
rect 420805 347454 421125 347486
rect 420805 347218 420847 347454
rect 421083 347218 421125 347454
rect 420805 347134 421125 347218
rect 420805 346898 420847 347134
rect 421083 346898 421125 347134
rect 420805 346866 421125 346898
rect 442874 347454 443194 347486
rect 442874 347218 442916 347454
rect 443152 347218 443194 347454
rect 442874 347134 443194 347218
rect 442874 346898 442916 347134
rect 443152 346898 443194 347134
rect 442874 346866 443194 346898
rect 448805 347454 449125 347486
rect 448805 347218 448847 347454
rect 449083 347218 449125 347454
rect 448805 347134 449125 347218
rect 448805 346898 448847 347134
rect 449083 346898 449125 347134
rect 448805 346866 449125 346898
rect 470874 347454 471194 347486
rect 470874 347218 470916 347454
rect 471152 347218 471194 347454
rect 470874 347134 471194 347218
rect 470874 346898 470916 347134
rect 471152 346898 471194 347134
rect 470874 346866 471194 346898
rect 476805 347454 477125 347486
rect 476805 347218 476847 347454
rect 477083 347218 477125 347454
rect 476805 347134 477125 347218
rect 476805 346898 476847 347134
rect 477083 346898 477125 347134
rect 476805 346866 477125 346898
rect 498874 347454 499194 347486
rect 498874 347218 498916 347454
rect 499152 347218 499194 347454
rect 498874 347134 499194 347218
rect 498874 346898 498916 347134
rect 499152 346898 499194 347134
rect 498874 346866 499194 346898
rect 504805 347454 505125 347486
rect 504805 347218 504847 347454
rect 505083 347218 505125 347454
rect 504805 347134 505125 347218
rect 504805 346898 504847 347134
rect 505083 346898 505125 347134
rect 504805 346866 505125 346898
rect 526874 347454 527194 347486
rect 526874 347218 526916 347454
rect 527152 347218 527194 347454
rect 526874 347134 527194 347218
rect 526874 346898 526916 347134
rect 527152 346898 527194 347134
rect 526874 346866 527194 346898
rect 532805 347454 533125 347486
rect 532805 347218 532847 347454
rect 533083 347218 533125 347454
rect 532805 347134 533125 347218
rect 532805 346898 532847 347134
rect 533083 346898 533125 347134
rect 532805 346866 533125 346898
rect 554874 347454 555194 347486
rect 554874 347218 554916 347454
rect 555152 347218 555194 347454
rect 554874 347134 555194 347218
rect 554874 346898 554916 347134
rect 555152 346898 555194 347134
rect 554874 346866 555194 346898
rect 560805 347454 561125 347486
rect 560805 347218 560847 347454
rect 561083 347218 561125 347454
rect 560805 347134 561125 347218
rect 560805 346898 560847 347134
rect 561083 346898 561125 347134
rect 560805 346866 561125 346898
rect -2006 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 -1386 323829
rect -2006 323509 -1386 323593
rect -2006 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 -1386 323509
rect -2006 296829 -1386 323273
rect 19910 323829 20230 323861
rect 19910 323593 19952 323829
rect 20188 323593 20230 323829
rect 19910 323509 20230 323593
rect 19910 323273 19952 323509
rect 20188 323273 20230 323509
rect 19910 323241 20230 323273
rect 25840 323829 26160 323861
rect 25840 323593 25882 323829
rect 26118 323593 26160 323829
rect 25840 323509 26160 323593
rect 25840 323273 25882 323509
rect 26118 323273 26160 323509
rect 25840 323241 26160 323273
rect 31771 323829 32091 323861
rect 31771 323593 31813 323829
rect 32049 323593 32091 323829
rect 31771 323509 32091 323593
rect 31771 323273 31813 323509
rect 32049 323273 32091 323509
rect 31771 323241 32091 323273
rect 47910 323829 48230 323861
rect 47910 323593 47952 323829
rect 48188 323593 48230 323829
rect 47910 323509 48230 323593
rect 47910 323273 47952 323509
rect 48188 323273 48230 323509
rect 47910 323241 48230 323273
rect 53840 323829 54160 323861
rect 53840 323593 53882 323829
rect 54118 323593 54160 323829
rect 53840 323509 54160 323593
rect 53840 323273 53882 323509
rect 54118 323273 54160 323509
rect 53840 323241 54160 323273
rect 59771 323829 60091 323861
rect 59771 323593 59813 323829
rect 60049 323593 60091 323829
rect 59771 323509 60091 323593
rect 59771 323273 59813 323509
rect 60049 323273 60091 323509
rect 59771 323241 60091 323273
rect 75910 323829 76230 323861
rect 75910 323593 75952 323829
rect 76188 323593 76230 323829
rect 75910 323509 76230 323593
rect 75910 323273 75952 323509
rect 76188 323273 76230 323509
rect 75910 323241 76230 323273
rect 81840 323829 82160 323861
rect 81840 323593 81882 323829
rect 82118 323593 82160 323829
rect 81840 323509 82160 323593
rect 81840 323273 81882 323509
rect 82118 323273 82160 323509
rect 81840 323241 82160 323273
rect 87771 323829 88091 323861
rect 87771 323593 87813 323829
rect 88049 323593 88091 323829
rect 87771 323509 88091 323593
rect 87771 323273 87813 323509
rect 88049 323273 88091 323509
rect 87771 323241 88091 323273
rect 103910 323829 104230 323861
rect 103910 323593 103952 323829
rect 104188 323593 104230 323829
rect 103910 323509 104230 323593
rect 103910 323273 103952 323509
rect 104188 323273 104230 323509
rect 103910 323241 104230 323273
rect 109840 323829 110160 323861
rect 109840 323593 109882 323829
rect 110118 323593 110160 323829
rect 109840 323509 110160 323593
rect 109840 323273 109882 323509
rect 110118 323273 110160 323509
rect 109840 323241 110160 323273
rect 115771 323829 116091 323861
rect 115771 323593 115813 323829
rect 116049 323593 116091 323829
rect 115771 323509 116091 323593
rect 115771 323273 115813 323509
rect 116049 323273 116091 323509
rect 115771 323241 116091 323273
rect 131910 323829 132230 323861
rect 131910 323593 131952 323829
rect 132188 323593 132230 323829
rect 131910 323509 132230 323593
rect 131910 323273 131952 323509
rect 132188 323273 132230 323509
rect 131910 323241 132230 323273
rect 137840 323829 138160 323861
rect 137840 323593 137882 323829
rect 138118 323593 138160 323829
rect 137840 323509 138160 323593
rect 137840 323273 137882 323509
rect 138118 323273 138160 323509
rect 137840 323241 138160 323273
rect 143771 323829 144091 323861
rect 143771 323593 143813 323829
rect 144049 323593 144091 323829
rect 143771 323509 144091 323593
rect 143771 323273 143813 323509
rect 144049 323273 144091 323509
rect 143771 323241 144091 323273
rect 159910 323829 160230 323861
rect 159910 323593 159952 323829
rect 160188 323593 160230 323829
rect 159910 323509 160230 323593
rect 159910 323273 159952 323509
rect 160188 323273 160230 323509
rect 159910 323241 160230 323273
rect 165840 323829 166160 323861
rect 165840 323593 165882 323829
rect 166118 323593 166160 323829
rect 165840 323509 166160 323593
rect 165840 323273 165882 323509
rect 166118 323273 166160 323509
rect 165840 323241 166160 323273
rect 171771 323829 172091 323861
rect 171771 323593 171813 323829
rect 172049 323593 172091 323829
rect 171771 323509 172091 323593
rect 171771 323273 171813 323509
rect 172049 323273 172091 323509
rect 171771 323241 172091 323273
rect 187910 323829 188230 323861
rect 187910 323593 187952 323829
rect 188188 323593 188230 323829
rect 187910 323509 188230 323593
rect 187910 323273 187952 323509
rect 188188 323273 188230 323509
rect 187910 323241 188230 323273
rect 193840 323829 194160 323861
rect 193840 323593 193882 323829
rect 194118 323593 194160 323829
rect 193840 323509 194160 323593
rect 193840 323273 193882 323509
rect 194118 323273 194160 323509
rect 193840 323241 194160 323273
rect 199771 323829 200091 323861
rect 199771 323593 199813 323829
rect 200049 323593 200091 323829
rect 199771 323509 200091 323593
rect 199771 323273 199813 323509
rect 200049 323273 200091 323509
rect 199771 323241 200091 323273
rect 215910 323829 216230 323861
rect 215910 323593 215952 323829
rect 216188 323593 216230 323829
rect 215910 323509 216230 323593
rect 215910 323273 215952 323509
rect 216188 323273 216230 323509
rect 215910 323241 216230 323273
rect 221840 323829 222160 323861
rect 221840 323593 221882 323829
rect 222118 323593 222160 323829
rect 221840 323509 222160 323593
rect 221840 323273 221882 323509
rect 222118 323273 222160 323509
rect 221840 323241 222160 323273
rect 227771 323829 228091 323861
rect 227771 323593 227813 323829
rect 228049 323593 228091 323829
rect 227771 323509 228091 323593
rect 227771 323273 227813 323509
rect 228049 323273 228091 323509
rect 227771 323241 228091 323273
rect 243910 323829 244230 323861
rect 243910 323593 243952 323829
rect 244188 323593 244230 323829
rect 243910 323509 244230 323593
rect 243910 323273 243952 323509
rect 244188 323273 244230 323509
rect 243910 323241 244230 323273
rect 249840 323829 250160 323861
rect 249840 323593 249882 323829
rect 250118 323593 250160 323829
rect 249840 323509 250160 323593
rect 249840 323273 249882 323509
rect 250118 323273 250160 323509
rect 249840 323241 250160 323273
rect 255771 323829 256091 323861
rect 255771 323593 255813 323829
rect 256049 323593 256091 323829
rect 255771 323509 256091 323593
rect 255771 323273 255813 323509
rect 256049 323273 256091 323509
rect 255771 323241 256091 323273
rect 271910 323829 272230 323861
rect 271910 323593 271952 323829
rect 272188 323593 272230 323829
rect 271910 323509 272230 323593
rect 271910 323273 271952 323509
rect 272188 323273 272230 323509
rect 271910 323241 272230 323273
rect 277840 323829 278160 323861
rect 277840 323593 277882 323829
rect 278118 323593 278160 323829
rect 277840 323509 278160 323593
rect 277840 323273 277882 323509
rect 278118 323273 278160 323509
rect 277840 323241 278160 323273
rect 283771 323829 284091 323861
rect 283771 323593 283813 323829
rect 284049 323593 284091 323829
rect 283771 323509 284091 323593
rect 283771 323273 283813 323509
rect 284049 323273 284091 323509
rect 283771 323241 284091 323273
rect 299910 323829 300230 323861
rect 299910 323593 299952 323829
rect 300188 323593 300230 323829
rect 299910 323509 300230 323593
rect 299910 323273 299952 323509
rect 300188 323273 300230 323509
rect 299910 323241 300230 323273
rect 305840 323829 306160 323861
rect 305840 323593 305882 323829
rect 306118 323593 306160 323829
rect 305840 323509 306160 323593
rect 305840 323273 305882 323509
rect 306118 323273 306160 323509
rect 305840 323241 306160 323273
rect 311771 323829 312091 323861
rect 311771 323593 311813 323829
rect 312049 323593 312091 323829
rect 311771 323509 312091 323593
rect 311771 323273 311813 323509
rect 312049 323273 312091 323509
rect 311771 323241 312091 323273
rect 327910 323829 328230 323861
rect 327910 323593 327952 323829
rect 328188 323593 328230 323829
rect 327910 323509 328230 323593
rect 327910 323273 327952 323509
rect 328188 323273 328230 323509
rect 327910 323241 328230 323273
rect 333840 323829 334160 323861
rect 333840 323593 333882 323829
rect 334118 323593 334160 323829
rect 333840 323509 334160 323593
rect 333840 323273 333882 323509
rect 334118 323273 334160 323509
rect 333840 323241 334160 323273
rect 339771 323829 340091 323861
rect 339771 323593 339813 323829
rect 340049 323593 340091 323829
rect 339771 323509 340091 323593
rect 339771 323273 339813 323509
rect 340049 323273 340091 323509
rect 339771 323241 340091 323273
rect 355910 323829 356230 323861
rect 355910 323593 355952 323829
rect 356188 323593 356230 323829
rect 355910 323509 356230 323593
rect 355910 323273 355952 323509
rect 356188 323273 356230 323509
rect 355910 323241 356230 323273
rect 361840 323829 362160 323861
rect 361840 323593 361882 323829
rect 362118 323593 362160 323829
rect 361840 323509 362160 323593
rect 361840 323273 361882 323509
rect 362118 323273 362160 323509
rect 361840 323241 362160 323273
rect 367771 323829 368091 323861
rect 367771 323593 367813 323829
rect 368049 323593 368091 323829
rect 367771 323509 368091 323593
rect 367771 323273 367813 323509
rect 368049 323273 368091 323509
rect 367771 323241 368091 323273
rect 383910 323829 384230 323861
rect 383910 323593 383952 323829
rect 384188 323593 384230 323829
rect 383910 323509 384230 323593
rect 383910 323273 383952 323509
rect 384188 323273 384230 323509
rect 383910 323241 384230 323273
rect 389840 323829 390160 323861
rect 389840 323593 389882 323829
rect 390118 323593 390160 323829
rect 389840 323509 390160 323593
rect 389840 323273 389882 323509
rect 390118 323273 390160 323509
rect 389840 323241 390160 323273
rect 395771 323829 396091 323861
rect 395771 323593 395813 323829
rect 396049 323593 396091 323829
rect 395771 323509 396091 323593
rect 395771 323273 395813 323509
rect 396049 323273 396091 323509
rect 395771 323241 396091 323273
rect 411910 323829 412230 323861
rect 411910 323593 411952 323829
rect 412188 323593 412230 323829
rect 411910 323509 412230 323593
rect 411910 323273 411952 323509
rect 412188 323273 412230 323509
rect 411910 323241 412230 323273
rect 417840 323829 418160 323861
rect 417840 323593 417882 323829
rect 418118 323593 418160 323829
rect 417840 323509 418160 323593
rect 417840 323273 417882 323509
rect 418118 323273 418160 323509
rect 417840 323241 418160 323273
rect 423771 323829 424091 323861
rect 423771 323593 423813 323829
rect 424049 323593 424091 323829
rect 423771 323509 424091 323593
rect 423771 323273 423813 323509
rect 424049 323273 424091 323509
rect 423771 323241 424091 323273
rect 439910 323829 440230 323861
rect 439910 323593 439952 323829
rect 440188 323593 440230 323829
rect 439910 323509 440230 323593
rect 439910 323273 439952 323509
rect 440188 323273 440230 323509
rect 439910 323241 440230 323273
rect 445840 323829 446160 323861
rect 445840 323593 445882 323829
rect 446118 323593 446160 323829
rect 445840 323509 446160 323593
rect 445840 323273 445882 323509
rect 446118 323273 446160 323509
rect 445840 323241 446160 323273
rect 451771 323829 452091 323861
rect 451771 323593 451813 323829
rect 452049 323593 452091 323829
rect 451771 323509 452091 323593
rect 451771 323273 451813 323509
rect 452049 323273 452091 323509
rect 451771 323241 452091 323273
rect 467910 323829 468230 323861
rect 467910 323593 467952 323829
rect 468188 323593 468230 323829
rect 467910 323509 468230 323593
rect 467910 323273 467952 323509
rect 468188 323273 468230 323509
rect 467910 323241 468230 323273
rect 473840 323829 474160 323861
rect 473840 323593 473882 323829
rect 474118 323593 474160 323829
rect 473840 323509 474160 323593
rect 473840 323273 473882 323509
rect 474118 323273 474160 323509
rect 473840 323241 474160 323273
rect 479771 323829 480091 323861
rect 479771 323593 479813 323829
rect 480049 323593 480091 323829
rect 479771 323509 480091 323593
rect 479771 323273 479813 323509
rect 480049 323273 480091 323509
rect 479771 323241 480091 323273
rect 495910 323829 496230 323861
rect 495910 323593 495952 323829
rect 496188 323593 496230 323829
rect 495910 323509 496230 323593
rect 495910 323273 495952 323509
rect 496188 323273 496230 323509
rect 495910 323241 496230 323273
rect 501840 323829 502160 323861
rect 501840 323593 501882 323829
rect 502118 323593 502160 323829
rect 501840 323509 502160 323593
rect 501840 323273 501882 323509
rect 502118 323273 502160 323509
rect 501840 323241 502160 323273
rect 507771 323829 508091 323861
rect 507771 323593 507813 323829
rect 508049 323593 508091 323829
rect 507771 323509 508091 323593
rect 507771 323273 507813 323509
rect 508049 323273 508091 323509
rect 507771 323241 508091 323273
rect 523910 323829 524230 323861
rect 523910 323593 523952 323829
rect 524188 323593 524230 323829
rect 523910 323509 524230 323593
rect 523910 323273 523952 323509
rect 524188 323273 524230 323509
rect 523910 323241 524230 323273
rect 529840 323829 530160 323861
rect 529840 323593 529882 323829
rect 530118 323593 530160 323829
rect 529840 323509 530160 323593
rect 529840 323273 529882 323509
rect 530118 323273 530160 323509
rect 529840 323241 530160 323273
rect 535771 323829 536091 323861
rect 535771 323593 535813 323829
rect 536049 323593 536091 323829
rect 535771 323509 536091 323593
rect 535771 323273 535813 323509
rect 536049 323273 536091 323509
rect 535771 323241 536091 323273
rect 551910 323829 552230 323861
rect 551910 323593 551952 323829
rect 552188 323593 552230 323829
rect 551910 323509 552230 323593
rect 551910 323273 551952 323509
rect 552188 323273 552230 323509
rect 551910 323241 552230 323273
rect 557840 323829 558160 323861
rect 557840 323593 557882 323829
rect 558118 323593 558160 323829
rect 557840 323509 558160 323593
rect 557840 323273 557882 323509
rect 558118 323273 558160 323509
rect 557840 323241 558160 323273
rect 563771 323829 564091 323861
rect 563771 323593 563813 323829
rect 564049 323593 564091 323829
rect 563771 323509 564091 323593
rect 563771 323273 563813 323509
rect 564049 323273 564091 323509
rect 563771 323241 564091 323273
rect 573494 323829 574114 350273
rect 573494 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 574114 323829
rect 573494 323509 574114 323593
rect 573494 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 574114 323509
rect 22874 320454 23194 320486
rect 22874 320218 22916 320454
rect 23152 320218 23194 320454
rect 22874 320134 23194 320218
rect 22874 319898 22916 320134
rect 23152 319898 23194 320134
rect 22874 319866 23194 319898
rect 28805 320454 29125 320486
rect 28805 320218 28847 320454
rect 29083 320218 29125 320454
rect 28805 320134 29125 320218
rect 28805 319898 28847 320134
rect 29083 319898 29125 320134
rect 28805 319866 29125 319898
rect 50874 320454 51194 320486
rect 50874 320218 50916 320454
rect 51152 320218 51194 320454
rect 50874 320134 51194 320218
rect 50874 319898 50916 320134
rect 51152 319898 51194 320134
rect 50874 319866 51194 319898
rect 56805 320454 57125 320486
rect 56805 320218 56847 320454
rect 57083 320218 57125 320454
rect 56805 320134 57125 320218
rect 56805 319898 56847 320134
rect 57083 319898 57125 320134
rect 56805 319866 57125 319898
rect 78874 320454 79194 320486
rect 78874 320218 78916 320454
rect 79152 320218 79194 320454
rect 78874 320134 79194 320218
rect 78874 319898 78916 320134
rect 79152 319898 79194 320134
rect 78874 319866 79194 319898
rect 84805 320454 85125 320486
rect 84805 320218 84847 320454
rect 85083 320218 85125 320454
rect 84805 320134 85125 320218
rect 84805 319898 84847 320134
rect 85083 319898 85125 320134
rect 84805 319866 85125 319898
rect 106874 320454 107194 320486
rect 106874 320218 106916 320454
rect 107152 320218 107194 320454
rect 106874 320134 107194 320218
rect 106874 319898 106916 320134
rect 107152 319898 107194 320134
rect 106874 319866 107194 319898
rect 112805 320454 113125 320486
rect 112805 320218 112847 320454
rect 113083 320218 113125 320454
rect 112805 320134 113125 320218
rect 112805 319898 112847 320134
rect 113083 319898 113125 320134
rect 112805 319866 113125 319898
rect 134874 320454 135194 320486
rect 134874 320218 134916 320454
rect 135152 320218 135194 320454
rect 134874 320134 135194 320218
rect 134874 319898 134916 320134
rect 135152 319898 135194 320134
rect 134874 319866 135194 319898
rect 140805 320454 141125 320486
rect 140805 320218 140847 320454
rect 141083 320218 141125 320454
rect 140805 320134 141125 320218
rect 140805 319898 140847 320134
rect 141083 319898 141125 320134
rect 140805 319866 141125 319898
rect 162874 320454 163194 320486
rect 162874 320218 162916 320454
rect 163152 320218 163194 320454
rect 162874 320134 163194 320218
rect 162874 319898 162916 320134
rect 163152 319898 163194 320134
rect 162874 319866 163194 319898
rect 168805 320454 169125 320486
rect 168805 320218 168847 320454
rect 169083 320218 169125 320454
rect 168805 320134 169125 320218
rect 168805 319898 168847 320134
rect 169083 319898 169125 320134
rect 168805 319866 169125 319898
rect 190874 320454 191194 320486
rect 190874 320218 190916 320454
rect 191152 320218 191194 320454
rect 190874 320134 191194 320218
rect 190874 319898 190916 320134
rect 191152 319898 191194 320134
rect 190874 319866 191194 319898
rect 196805 320454 197125 320486
rect 196805 320218 196847 320454
rect 197083 320218 197125 320454
rect 196805 320134 197125 320218
rect 196805 319898 196847 320134
rect 197083 319898 197125 320134
rect 196805 319866 197125 319898
rect 218874 320454 219194 320486
rect 218874 320218 218916 320454
rect 219152 320218 219194 320454
rect 218874 320134 219194 320218
rect 218874 319898 218916 320134
rect 219152 319898 219194 320134
rect 218874 319866 219194 319898
rect 224805 320454 225125 320486
rect 224805 320218 224847 320454
rect 225083 320218 225125 320454
rect 224805 320134 225125 320218
rect 224805 319898 224847 320134
rect 225083 319898 225125 320134
rect 224805 319866 225125 319898
rect 246874 320454 247194 320486
rect 246874 320218 246916 320454
rect 247152 320218 247194 320454
rect 246874 320134 247194 320218
rect 246874 319898 246916 320134
rect 247152 319898 247194 320134
rect 246874 319866 247194 319898
rect 252805 320454 253125 320486
rect 252805 320218 252847 320454
rect 253083 320218 253125 320454
rect 252805 320134 253125 320218
rect 252805 319898 252847 320134
rect 253083 319898 253125 320134
rect 252805 319866 253125 319898
rect 274874 320454 275194 320486
rect 274874 320218 274916 320454
rect 275152 320218 275194 320454
rect 274874 320134 275194 320218
rect 274874 319898 274916 320134
rect 275152 319898 275194 320134
rect 274874 319866 275194 319898
rect 280805 320454 281125 320486
rect 280805 320218 280847 320454
rect 281083 320218 281125 320454
rect 280805 320134 281125 320218
rect 280805 319898 280847 320134
rect 281083 319898 281125 320134
rect 280805 319866 281125 319898
rect 302874 320454 303194 320486
rect 302874 320218 302916 320454
rect 303152 320218 303194 320454
rect 302874 320134 303194 320218
rect 302874 319898 302916 320134
rect 303152 319898 303194 320134
rect 302874 319866 303194 319898
rect 308805 320454 309125 320486
rect 308805 320218 308847 320454
rect 309083 320218 309125 320454
rect 308805 320134 309125 320218
rect 308805 319898 308847 320134
rect 309083 319898 309125 320134
rect 308805 319866 309125 319898
rect 330874 320454 331194 320486
rect 330874 320218 330916 320454
rect 331152 320218 331194 320454
rect 330874 320134 331194 320218
rect 330874 319898 330916 320134
rect 331152 319898 331194 320134
rect 330874 319866 331194 319898
rect 336805 320454 337125 320486
rect 336805 320218 336847 320454
rect 337083 320218 337125 320454
rect 336805 320134 337125 320218
rect 336805 319898 336847 320134
rect 337083 319898 337125 320134
rect 336805 319866 337125 319898
rect 358874 320454 359194 320486
rect 358874 320218 358916 320454
rect 359152 320218 359194 320454
rect 358874 320134 359194 320218
rect 358874 319898 358916 320134
rect 359152 319898 359194 320134
rect 358874 319866 359194 319898
rect 364805 320454 365125 320486
rect 364805 320218 364847 320454
rect 365083 320218 365125 320454
rect 364805 320134 365125 320218
rect 364805 319898 364847 320134
rect 365083 319898 365125 320134
rect 364805 319866 365125 319898
rect 386874 320454 387194 320486
rect 386874 320218 386916 320454
rect 387152 320218 387194 320454
rect 386874 320134 387194 320218
rect 386874 319898 386916 320134
rect 387152 319898 387194 320134
rect 386874 319866 387194 319898
rect 392805 320454 393125 320486
rect 392805 320218 392847 320454
rect 393083 320218 393125 320454
rect 392805 320134 393125 320218
rect 392805 319898 392847 320134
rect 393083 319898 393125 320134
rect 392805 319866 393125 319898
rect 414874 320454 415194 320486
rect 414874 320218 414916 320454
rect 415152 320218 415194 320454
rect 414874 320134 415194 320218
rect 414874 319898 414916 320134
rect 415152 319898 415194 320134
rect 414874 319866 415194 319898
rect 420805 320454 421125 320486
rect 420805 320218 420847 320454
rect 421083 320218 421125 320454
rect 420805 320134 421125 320218
rect 420805 319898 420847 320134
rect 421083 319898 421125 320134
rect 420805 319866 421125 319898
rect 442874 320454 443194 320486
rect 442874 320218 442916 320454
rect 443152 320218 443194 320454
rect 442874 320134 443194 320218
rect 442874 319898 442916 320134
rect 443152 319898 443194 320134
rect 442874 319866 443194 319898
rect 448805 320454 449125 320486
rect 448805 320218 448847 320454
rect 449083 320218 449125 320454
rect 448805 320134 449125 320218
rect 448805 319898 448847 320134
rect 449083 319898 449125 320134
rect 448805 319866 449125 319898
rect 470874 320454 471194 320486
rect 470874 320218 470916 320454
rect 471152 320218 471194 320454
rect 470874 320134 471194 320218
rect 470874 319898 470916 320134
rect 471152 319898 471194 320134
rect 470874 319866 471194 319898
rect 476805 320454 477125 320486
rect 476805 320218 476847 320454
rect 477083 320218 477125 320454
rect 476805 320134 477125 320218
rect 476805 319898 476847 320134
rect 477083 319898 477125 320134
rect 476805 319866 477125 319898
rect 498874 320454 499194 320486
rect 498874 320218 498916 320454
rect 499152 320218 499194 320454
rect 498874 320134 499194 320218
rect 498874 319898 498916 320134
rect 499152 319898 499194 320134
rect 498874 319866 499194 319898
rect 504805 320454 505125 320486
rect 504805 320218 504847 320454
rect 505083 320218 505125 320454
rect 504805 320134 505125 320218
rect 504805 319898 504847 320134
rect 505083 319898 505125 320134
rect 504805 319866 505125 319898
rect 526874 320454 527194 320486
rect 526874 320218 526916 320454
rect 527152 320218 527194 320454
rect 526874 320134 527194 320218
rect 526874 319898 526916 320134
rect 527152 319898 527194 320134
rect 526874 319866 527194 319898
rect 532805 320454 533125 320486
rect 532805 320218 532847 320454
rect 533083 320218 533125 320454
rect 532805 320134 533125 320218
rect 532805 319898 532847 320134
rect 533083 319898 533125 320134
rect 532805 319866 533125 319898
rect 554874 320454 555194 320486
rect 554874 320218 554916 320454
rect 555152 320218 555194 320454
rect 554874 320134 555194 320218
rect 554874 319898 554916 320134
rect 555152 319898 555194 320134
rect 554874 319866 555194 319898
rect 560805 320454 561125 320486
rect 560805 320218 560847 320454
rect 561083 320218 561125 320454
rect 560805 320134 561125 320218
rect 560805 319898 560847 320134
rect 561083 319898 561125 320134
rect 560805 319866 561125 319898
rect -2006 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 -1386 296829
rect -2006 296509 -1386 296593
rect -2006 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 -1386 296509
rect -2006 269829 -1386 296273
rect 19910 296829 20230 296861
rect 19910 296593 19952 296829
rect 20188 296593 20230 296829
rect 19910 296509 20230 296593
rect 19910 296273 19952 296509
rect 20188 296273 20230 296509
rect 19910 296241 20230 296273
rect 25840 296829 26160 296861
rect 25840 296593 25882 296829
rect 26118 296593 26160 296829
rect 25840 296509 26160 296593
rect 25840 296273 25882 296509
rect 26118 296273 26160 296509
rect 25840 296241 26160 296273
rect 31771 296829 32091 296861
rect 31771 296593 31813 296829
rect 32049 296593 32091 296829
rect 31771 296509 32091 296593
rect 31771 296273 31813 296509
rect 32049 296273 32091 296509
rect 31771 296241 32091 296273
rect 47910 296829 48230 296861
rect 47910 296593 47952 296829
rect 48188 296593 48230 296829
rect 47910 296509 48230 296593
rect 47910 296273 47952 296509
rect 48188 296273 48230 296509
rect 47910 296241 48230 296273
rect 53840 296829 54160 296861
rect 53840 296593 53882 296829
rect 54118 296593 54160 296829
rect 53840 296509 54160 296593
rect 53840 296273 53882 296509
rect 54118 296273 54160 296509
rect 53840 296241 54160 296273
rect 59771 296829 60091 296861
rect 59771 296593 59813 296829
rect 60049 296593 60091 296829
rect 59771 296509 60091 296593
rect 59771 296273 59813 296509
rect 60049 296273 60091 296509
rect 59771 296241 60091 296273
rect 75910 296829 76230 296861
rect 75910 296593 75952 296829
rect 76188 296593 76230 296829
rect 75910 296509 76230 296593
rect 75910 296273 75952 296509
rect 76188 296273 76230 296509
rect 75910 296241 76230 296273
rect 81840 296829 82160 296861
rect 81840 296593 81882 296829
rect 82118 296593 82160 296829
rect 81840 296509 82160 296593
rect 81840 296273 81882 296509
rect 82118 296273 82160 296509
rect 81840 296241 82160 296273
rect 87771 296829 88091 296861
rect 87771 296593 87813 296829
rect 88049 296593 88091 296829
rect 87771 296509 88091 296593
rect 87771 296273 87813 296509
rect 88049 296273 88091 296509
rect 87771 296241 88091 296273
rect 103910 296829 104230 296861
rect 103910 296593 103952 296829
rect 104188 296593 104230 296829
rect 103910 296509 104230 296593
rect 103910 296273 103952 296509
rect 104188 296273 104230 296509
rect 103910 296241 104230 296273
rect 109840 296829 110160 296861
rect 109840 296593 109882 296829
rect 110118 296593 110160 296829
rect 109840 296509 110160 296593
rect 109840 296273 109882 296509
rect 110118 296273 110160 296509
rect 109840 296241 110160 296273
rect 115771 296829 116091 296861
rect 115771 296593 115813 296829
rect 116049 296593 116091 296829
rect 115771 296509 116091 296593
rect 115771 296273 115813 296509
rect 116049 296273 116091 296509
rect 115771 296241 116091 296273
rect 131910 296829 132230 296861
rect 131910 296593 131952 296829
rect 132188 296593 132230 296829
rect 131910 296509 132230 296593
rect 131910 296273 131952 296509
rect 132188 296273 132230 296509
rect 131910 296241 132230 296273
rect 137840 296829 138160 296861
rect 137840 296593 137882 296829
rect 138118 296593 138160 296829
rect 137840 296509 138160 296593
rect 137840 296273 137882 296509
rect 138118 296273 138160 296509
rect 137840 296241 138160 296273
rect 143771 296829 144091 296861
rect 143771 296593 143813 296829
rect 144049 296593 144091 296829
rect 143771 296509 144091 296593
rect 143771 296273 143813 296509
rect 144049 296273 144091 296509
rect 143771 296241 144091 296273
rect 159910 296829 160230 296861
rect 159910 296593 159952 296829
rect 160188 296593 160230 296829
rect 159910 296509 160230 296593
rect 159910 296273 159952 296509
rect 160188 296273 160230 296509
rect 159910 296241 160230 296273
rect 165840 296829 166160 296861
rect 165840 296593 165882 296829
rect 166118 296593 166160 296829
rect 165840 296509 166160 296593
rect 165840 296273 165882 296509
rect 166118 296273 166160 296509
rect 165840 296241 166160 296273
rect 171771 296829 172091 296861
rect 171771 296593 171813 296829
rect 172049 296593 172091 296829
rect 171771 296509 172091 296593
rect 171771 296273 171813 296509
rect 172049 296273 172091 296509
rect 171771 296241 172091 296273
rect 187910 296829 188230 296861
rect 187910 296593 187952 296829
rect 188188 296593 188230 296829
rect 187910 296509 188230 296593
rect 187910 296273 187952 296509
rect 188188 296273 188230 296509
rect 187910 296241 188230 296273
rect 193840 296829 194160 296861
rect 193840 296593 193882 296829
rect 194118 296593 194160 296829
rect 193840 296509 194160 296593
rect 193840 296273 193882 296509
rect 194118 296273 194160 296509
rect 193840 296241 194160 296273
rect 199771 296829 200091 296861
rect 199771 296593 199813 296829
rect 200049 296593 200091 296829
rect 199771 296509 200091 296593
rect 199771 296273 199813 296509
rect 200049 296273 200091 296509
rect 199771 296241 200091 296273
rect 215910 296829 216230 296861
rect 215910 296593 215952 296829
rect 216188 296593 216230 296829
rect 215910 296509 216230 296593
rect 215910 296273 215952 296509
rect 216188 296273 216230 296509
rect 215910 296241 216230 296273
rect 221840 296829 222160 296861
rect 221840 296593 221882 296829
rect 222118 296593 222160 296829
rect 221840 296509 222160 296593
rect 221840 296273 221882 296509
rect 222118 296273 222160 296509
rect 221840 296241 222160 296273
rect 227771 296829 228091 296861
rect 227771 296593 227813 296829
rect 228049 296593 228091 296829
rect 227771 296509 228091 296593
rect 227771 296273 227813 296509
rect 228049 296273 228091 296509
rect 227771 296241 228091 296273
rect 243910 296829 244230 296861
rect 243910 296593 243952 296829
rect 244188 296593 244230 296829
rect 243910 296509 244230 296593
rect 243910 296273 243952 296509
rect 244188 296273 244230 296509
rect 243910 296241 244230 296273
rect 249840 296829 250160 296861
rect 249840 296593 249882 296829
rect 250118 296593 250160 296829
rect 249840 296509 250160 296593
rect 249840 296273 249882 296509
rect 250118 296273 250160 296509
rect 249840 296241 250160 296273
rect 255771 296829 256091 296861
rect 255771 296593 255813 296829
rect 256049 296593 256091 296829
rect 255771 296509 256091 296593
rect 255771 296273 255813 296509
rect 256049 296273 256091 296509
rect 255771 296241 256091 296273
rect 271910 296829 272230 296861
rect 271910 296593 271952 296829
rect 272188 296593 272230 296829
rect 271910 296509 272230 296593
rect 271910 296273 271952 296509
rect 272188 296273 272230 296509
rect 271910 296241 272230 296273
rect 277840 296829 278160 296861
rect 277840 296593 277882 296829
rect 278118 296593 278160 296829
rect 277840 296509 278160 296593
rect 277840 296273 277882 296509
rect 278118 296273 278160 296509
rect 277840 296241 278160 296273
rect 283771 296829 284091 296861
rect 283771 296593 283813 296829
rect 284049 296593 284091 296829
rect 283771 296509 284091 296593
rect 283771 296273 283813 296509
rect 284049 296273 284091 296509
rect 283771 296241 284091 296273
rect 299910 296829 300230 296861
rect 299910 296593 299952 296829
rect 300188 296593 300230 296829
rect 299910 296509 300230 296593
rect 299910 296273 299952 296509
rect 300188 296273 300230 296509
rect 299910 296241 300230 296273
rect 305840 296829 306160 296861
rect 305840 296593 305882 296829
rect 306118 296593 306160 296829
rect 305840 296509 306160 296593
rect 305840 296273 305882 296509
rect 306118 296273 306160 296509
rect 305840 296241 306160 296273
rect 311771 296829 312091 296861
rect 311771 296593 311813 296829
rect 312049 296593 312091 296829
rect 311771 296509 312091 296593
rect 311771 296273 311813 296509
rect 312049 296273 312091 296509
rect 311771 296241 312091 296273
rect 327910 296829 328230 296861
rect 327910 296593 327952 296829
rect 328188 296593 328230 296829
rect 327910 296509 328230 296593
rect 327910 296273 327952 296509
rect 328188 296273 328230 296509
rect 327910 296241 328230 296273
rect 333840 296829 334160 296861
rect 333840 296593 333882 296829
rect 334118 296593 334160 296829
rect 333840 296509 334160 296593
rect 333840 296273 333882 296509
rect 334118 296273 334160 296509
rect 333840 296241 334160 296273
rect 339771 296829 340091 296861
rect 339771 296593 339813 296829
rect 340049 296593 340091 296829
rect 339771 296509 340091 296593
rect 339771 296273 339813 296509
rect 340049 296273 340091 296509
rect 339771 296241 340091 296273
rect 355910 296829 356230 296861
rect 355910 296593 355952 296829
rect 356188 296593 356230 296829
rect 355910 296509 356230 296593
rect 355910 296273 355952 296509
rect 356188 296273 356230 296509
rect 355910 296241 356230 296273
rect 361840 296829 362160 296861
rect 361840 296593 361882 296829
rect 362118 296593 362160 296829
rect 361840 296509 362160 296593
rect 361840 296273 361882 296509
rect 362118 296273 362160 296509
rect 361840 296241 362160 296273
rect 367771 296829 368091 296861
rect 367771 296593 367813 296829
rect 368049 296593 368091 296829
rect 367771 296509 368091 296593
rect 367771 296273 367813 296509
rect 368049 296273 368091 296509
rect 367771 296241 368091 296273
rect 383910 296829 384230 296861
rect 383910 296593 383952 296829
rect 384188 296593 384230 296829
rect 383910 296509 384230 296593
rect 383910 296273 383952 296509
rect 384188 296273 384230 296509
rect 383910 296241 384230 296273
rect 389840 296829 390160 296861
rect 389840 296593 389882 296829
rect 390118 296593 390160 296829
rect 389840 296509 390160 296593
rect 389840 296273 389882 296509
rect 390118 296273 390160 296509
rect 389840 296241 390160 296273
rect 395771 296829 396091 296861
rect 395771 296593 395813 296829
rect 396049 296593 396091 296829
rect 395771 296509 396091 296593
rect 395771 296273 395813 296509
rect 396049 296273 396091 296509
rect 395771 296241 396091 296273
rect 411910 296829 412230 296861
rect 411910 296593 411952 296829
rect 412188 296593 412230 296829
rect 411910 296509 412230 296593
rect 411910 296273 411952 296509
rect 412188 296273 412230 296509
rect 411910 296241 412230 296273
rect 417840 296829 418160 296861
rect 417840 296593 417882 296829
rect 418118 296593 418160 296829
rect 417840 296509 418160 296593
rect 417840 296273 417882 296509
rect 418118 296273 418160 296509
rect 417840 296241 418160 296273
rect 423771 296829 424091 296861
rect 423771 296593 423813 296829
rect 424049 296593 424091 296829
rect 423771 296509 424091 296593
rect 423771 296273 423813 296509
rect 424049 296273 424091 296509
rect 423771 296241 424091 296273
rect 439910 296829 440230 296861
rect 439910 296593 439952 296829
rect 440188 296593 440230 296829
rect 439910 296509 440230 296593
rect 439910 296273 439952 296509
rect 440188 296273 440230 296509
rect 439910 296241 440230 296273
rect 445840 296829 446160 296861
rect 445840 296593 445882 296829
rect 446118 296593 446160 296829
rect 445840 296509 446160 296593
rect 445840 296273 445882 296509
rect 446118 296273 446160 296509
rect 445840 296241 446160 296273
rect 451771 296829 452091 296861
rect 451771 296593 451813 296829
rect 452049 296593 452091 296829
rect 451771 296509 452091 296593
rect 451771 296273 451813 296509
rect 452049 296273 452091 296509
rect 451771 296241 452091 296273
rect 467910 296829 468230 296861
rect 467910 296593 467952 296829
rect 468188 296593 468230 296829
rect 467910 296509 468230 296593
rect 467910 296273 467952 296509
rect 468188 296273 468230 296509
rect 467910 296241 468230 296273
rect 473840 296829 474160 296861
rect 473840 296593 473882 296829
rect 474118 296593 474160 296829
rect 473840 296509 474160 296593
rect 473840 296273 473882 296509
rect 474118 296273 474160 296509
rect 473840 296241 474160 296273
rect 479771 296829 480091 296861
rect 479771 296593 479813 296829
rect 480049 296593 480091 296829
rect 479771 296509 480091 296593
rect 479771 296273 479813 296509
rect 480049 296273 480091 296509
rect 479771 296241 480091 296273
rect 495910 296829 496230 296861
rect 495910 296593 495952 296829
rect 496188 296593 496230 296829
rect 495910 296509 496230 296593
rect 495910 296273 495952 296509
rect 496188 296273 496230 296509
rect 495910 296241 496230 296273
rect 501840 296829 502160 296861
rect 501840 296593 501882 296829
rect 502118 296593 502160 296829
rect 501840 296509 502160 296593
rect 501840 296273 501882 296509
rect 502118 296273 502160 296509
rect 501840 296241 502160 296273
rect 507771 296829 508091 296861
rect 507771 296593 507813 296829
rect 508049 296593 508091 296829
rect 507771 296509 508091 296593
rect 507771 296273 507813 296509
rect 508049 296273 508091 296509
rect 507771 296241 508091 296273
rect 523910 296829 524230 296861
rect 523910 296593 523952 296829
rect 524188 296593 524230 296829
rect 523910 296509 524230 296593
rect 523910 296273 523952 296509
rect 524188 296273 524230 296509
rect 523910 296241 524230 296273
rect 529840 296829 530160 296861
rect 529840 296593 529882 296829
rect 530118 296593 530160 296829
rect 529840 296509 530160 296593
rect 529840 296273 529882 296509
rect 530118 296273 530160 296509
rect 529840 296241 530160 296273
rect 535771 296829 536091 296861
rect 535771 296593 535813 296829
rect 536049 296593 536091 296829
rect 535771 296509 536091 296593
rect 535771 296273 535813 296509
rect 536049 296273 536091 296509
rect 535771 296241 536091 296273
rect 551910 296829 552230 296861
rect 551910 296593 551952 296829
rect 552188 296593 552230 296829
rect 551910 296509 552230 296593
rect 551910 296273 551952 296509
rect 552188 296273 552230 296509
rect 551910 296241 552230 296273
rect 557840 296829 558160 296861
rect 557840 296593 557882 296829
rect 558118 296593 558160 296829
rect 557840 296509 558160 296593
rect 557840 296273 557882 296509
rect 558118 296273 558160 296509
rect 557840 296241 558160 296273
rect 563771 296829 564091 296861
rect 563771 296593 563813 296829
rect 564049 296593 564091 296829
rect 563771 296509 564091 296593
rect 563771 296273 563813 296509
rect 564049 296273 564091 296509
rect 563771 296241 564091 296273
rect 573494 296829 574114 323273
rect 573494 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 574114 296829
rect 573494 296509 574114 296593
rect 573494 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 574114 296509
rect 22874 293454 23194 293486
rect 22874 293218 22916 293454
rect 23152 293218 23194 293454
rect 22874 293134 23194 293218
rect 22874 292898 22916 293134
rect 23152 292898 23194 293134
rect 22874 292866 23194 292898
rect 28805 293454 29125 293486
rect 28805 293218 28847 293454
rect 29083 293218 29125 293454
rect 28805 293134 29125 293218
rect 28805 292898 28847 293134
rect 29083 292898 29125 293134
rect 28805 292866 29125 292898
rect 50874 293454 51194 293486
rect 50874 293218 50916 293454
rect 51152 293218 51194 293454
rect 50874 293134 51194 293218
rect 50874 292898 50916 293134
rect 51152 292898 51194 293134
rect 50874 292866 51194 292898
rect 56805 293454 57125 293486
rect 56805 293218 56847 293454
rect 57083 293218 57125 293454
rect 56805 293134 57125 293218
rect 56805 292898 56847 293134
rect 57083 292898 57125 293134
rect 56805 292866 57125 292898
rect 78874 293454 79194 293486
rect 78874 293218 78916 293454
rect 79152 293218 79194 293454
rect 78874 293134 79194 293218
rect 78874 292898 78916 293134
rect 79152 292898 79194 293134
rect 78874 292866 79194 292898
rect 84805 293454 85125 293486
rect 84805 293218 84847 293454
rect 85083 293218 85125 293454
rect 84805 293134 85125 293218
rect 84805 292898 84847 293134
rect 85083 292898 85125 293134
rect 84805 292866 85125 292898
rect 106874 293454 107194 293486
rect 106874 293218 106916 293454
rect 107152 293218 107194 293454
rect 106874 293134 107194 293218
rect 106874 292898 106916 293134
rect 107152 292898 107194 293134
rect 106874 292866 107194 292898
rect 112805 293454 113125 293486
rect 112805 293218 112847 293454
rect 113083 293218 113125 293454
rect 112805 293134 113125 293218
rect 112805 292898 112847 293134
rect 113083 292898 113125 293134
rect 112805 292866 113125 292898
rect 134874 293454 135194 293486
rect 134874 293218 134916 293454
rect 135152 293218 135194 293454
rect 134874 293134 135194 293218
rect 134874 292898 134916 293134
rect 135152 292898 135194 293134
rect 134874 292866 135194 292898
rect 140805 293454 141125 293486
rect 140805 293218 140847 293454
rect 141083 293218 141125 293454
rect 140805 293134 141125 293218
rect 140805 292898 140847 293134
rect 141083 292898 141125 293134
rect 140805 292866 141125 292898
rect 162874 293454 163194 293486
rect 162874 293218 162916 293454
rect 163152 293218 163194 293454
rect 162874 293134 163194 293218
rect 162874 292898 162916 293134
rect 163152 292898 163194 293134
rect 162874 292866 163194 292898
rect 168805 293454 169125 293486
rect 168805 293218 168847 293454
rect 169083 293218 169125 293454
rect 168805 293134 169125 293218
rect 168805 292898 168847 293134
rect 169083 292898 169125 293134
rect 168805 292866 169125 292898
rect 190874 293454 191194 293486
rect 190874 293218 190916 293454
rect 191152 293218 191194 293454
rect 190874 293134 191194 293218
rect 190874 292898 190916 293134
rect 191152 292898 191194 293134
rect 190874 292866 191194 292898
rect 196805 293454 197125 293486
rect 196805 293218 196847 293454
rect 197083 293218 197125 293454
rect 196805 293134 197125 293218
rect 196805 292898 196847 293134
rect 197083 292898 197125 293134
rect 196805 292866 197125 292898
rect 218874 293454 219194 293486
rect 218874 293218 218916 293454
rect 219152 293218 219194 293454
rect 218874 293134 219194 293218
rect 218874 292898 218916 293134
rect 219152 292898 219194 293134
rect 218874 292866 219194 292898
rect 224805 293454 225125 293486
rect 224805 293218 224847 293454
rect 225083 293218 225125 293454
rect 224805 293134 225125 293218
rect 224805 292898 224847 293134
rect 225083 292898 225125 293134
rect 224805 292866 225125 292898
rect 246874 293454 247194 293486
rect 246874 293218 246916 293454
rect 247152 293218 247194 293454
rect 246874 293134 247194 293218
rect 246874 292898 246916 293134
rect 247152 292898 247194 293134
rect 246874 292866 247194 292898
rect 252805 293454 253125 293486
rect 252805 293218 252847 293454
rect 253083 293218 253125 293454
rect 252805 293134 253125 293218
rect 252805 292898 252847 293134
rect 253083 292898 253125 293134
rect 252805 292866 253125 292898
rect 274874 293454 275194 293486
rect 274874 293218 274916 293454
rect 275152 293218 275194 293454
rect 274874 293134 275194 293218
rect 274874 292898 274916 293134
rect 275152 292898 275194 293134
rect 274874 292866 275194 292898
rect 280805 293454 281125 293486
rect 280805 293218 280847 293454
rect 281083 293218 281125 293454
rect 280805 293134 281125 293218
rect 280805 292898 280847 293134
rect 281083 292898 281125 293134
rect 280805 292866 281125 292898
rect 302874 293454 303194 293486
rect 302874 293218 302916 293454
rect 303152 293218 303194 293454
rect 302874 293134 303194 293218
rect 302874 292898 302916 293134
rect 303152 292898 303194 293134
rect 302874 292866 303194 292898
rect 308805 293454 309125 293486
rect 308805 293218 308847 293454
rect 309083 293218 309125 293454
rect 308805 293134 309125 293218
rect 308805 292898 308847 293134
rect 309083 292898 309125 293134
rect 308805 292866 309125 292898
rect 330874 293454 331194 293486
rect 330874 293218 330916 293454
rect 331152 293218 331194 293454
rect 330874 293134 331194 293218
rect 330874 292898 330916 293134
rect 331152 292898 331194 293134
rect 330874 292866 331194 292898
rect 336805 293454 337125 293486
rect 336805 293218 336847 293454
rect 337083 293218 337125 293454
rect 336805 293134 337125 293218
rect 336805 292898 336847 293134
rect 337083 292898 337125 293134
rect 336805 292866 337125 292898
rect 358874 293454 359194 293486
rect 358874 293218 358916 293454
rect 359152 293218 359194 293454
rect 358874 293134 359194 293218
rect 358874 292898 358916 293134
rect 359152 292898 359194 293134
rect 358874 292866 359194 292898
rect 364805 293454 365125 293486
rect 364805 293218 364847 293454
rect 365083 293218 365125 293454
rect 364805 293134 365125 293218
rect 364805 292898 364847 293134
rect 365083 292898 365125 293134
rect 364805 292866 365125 292898
rect 386874 293454 387194 293486
rect 386874 293218 386916 293454
rect 387152 293218 387194 293454
rect 386874 293134 387194 293218
rect 386874 292898 386916 293134
rect 387152 292898 387194 293134
rect 386874 292866 387194 292898
rect 392805 293454 393125 293486
rect 392805 293218 392847 293454
rect 393083 293218 393125 293454
rect 392805 293134 393125 293218
rect 392805 292898 392847 293134
rect 393083 292898 393125 293134
rect 392805 292866 393125 292898
rect 414874 293454 415194 293486
rect 414874 293218 414916 293454
rect 415152 293218 415194 293454
rect 414874 293134 415194 293218
rect 414874 292898 414916 293134
rect 415152 292898 415194 293134
rect 414874 292866 415194 292898
rect 420805 293454 421125 293486
rect 420805 293218 420847 293454
rect 421083 293218 421125 293454
rect 420805 293134 421125 293218
rect 420805 292898 420847 293134
rect 421083 292898 421125 293134
rect 420805 292866 421125 292898
rect 442874 293454 443194 293486
rect 442874 293218 442916 293454
rect 443152 293218 443194 293454
rect 442874 293134 443194 293218
rect 442874 292898 442916 293134
rect 443152 292898 443194 293134
rect 442874 292866 443194 292898
rect 448805 293454 449125 293486
rect 448805 293218 448847 293454
rect 449083 293218 449125 293454
rect 448805 293134 449125 293218
rect 448805 292898 448847 293134
rect 449083 292898 449125 293134
rect 448805 292866 449125 292898
rect 470874 293454 471194 293486
rect 470874 293218 470916 293454
rect 471152 293218 471194 293454
rect 470874 293134 471194 293218
rect 470874 292898 470916 293134
rect 471152 292898 471194 293134
rect 470874 292866 471194 292898
rect 476805 293454 477125 293486
rect 476805 293218 476847 293454
rect 477083 293218 477125 293454
rect 476805 293134 477125 293218
rect 476805 292898 476847 293134
rect 477083 292898 477125 293134
rect 476805 292866 477125 292898
rect 498874 293454 499194 293486
rect 498874 293218 498916 293454
rect 499152 293218 499194 293454
rect 498874 293134 499194 293218
rect 498874 292898 498916 293134
rect 499152 292898 499194 293134
rect 498874 292866 499194 292898
rect 504805 293454 505125 293486
rect 504805 293218 504847 293454
rect 505083 293218 505125 293454
rect 504805 293134 505125 293218
rect 504805 292898 504847 293134
rect 505083 292898 505125 293134
rect 504805 292866 505125 292898
rect 526874 293454 527194 293486
rect 526874 293218 526916 293454
rect 527152 293218 527194 293454
rect 526874 293134 527194 293218
rect 526874 292898 526916 293134
rect 527152 292898 527194 293134
rect 526874 292866 527194 292898
rect 532805 293454 533125 293486
rect 532805 293218 532847 293454
rect 533083 293218 533125 293454
rect 532805 293134 533125 293218
rect 532805 292898 532847 293134
rect 533083 292898 533125 293134
rect 532805 292866 533125 292898
rect 554874 293454 555194 293486
rect 554874 293218 554916 293454
rect 555152 293218 555194 293454
rect 554874 293134 555194 293218
rect 554874 292898 554916 293134
rect 555152 292898 555194 293134
rect 554874 292866 555194 292898
rect 560805 293454 561125 293486
rect 560805 293218 560847 293454
rect 561083 293218 561125 293454
rect 560805 293134 561125 293218
rect 560805 292898 560847 293134
rect 561083 292898 561125 293134
rect 560805 292866 561125 292898
rect -2006 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 -1386 269829
rect -2006 269509 -1386 269593
rect -2006 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 -1386 269509
rect -2006 242829 -1386 269273
rect 19910 269829 20230 269861
rect 19910 269593 19952 269829
rect 20188 269593 20230 269829
rect 19910 269509 20230 269593
rect 19910 269273 19952 269509
rect 20188 269273 20230 269509
rect 19910 269241 20230 269273
rect 25840 269829 26160 269861
rect 25840 269593 25882 269829
rect 26118 269593 26160 269829
rect 25840 269509 26160 269593
rect 25840 269273 25882 269509
rect 26118 269273 26160 269509
rect 25840 269241 26160 269273
rect 31771 269829 32091 269861
rect 31771 269593 31813 269829
rect 32049 269593 32091 269829
rect 31771 269509 32091 269593
rect 31771 269273 31813 269509
rect 32049 269273 32091 269509
rect 31771 269241 32091 269273
rect 47910 269829 48230 269861
rect 47910 269593 47952 269829
rect 48188 269593 48230 269829
rect 47910 269509 48230 269593
rect 47910 269273 47952 269509
rect 48188 269273 48230 269509
rect 47910 269241 48230 269273
rect 53840 269829 54160 269861
rect 53840 269593 53882 269829
rect 54118 269593 54160 269829
rect 53840 269509 54160 269593
rect 53840 269273 53882 269509
rect 54118 269273 54160 269509
rect 53840 269241 54160 269273
rect 59771 269829 60091 269861
rect 59771 269593 59813 269829
rect 60049 269593 60091 269829
rect 59771 269509 60091 269593
rect 59771 269273 59813 269509
rect 60049 269273 60091 269509
rect 59771 269241 60091 269273
rect 75910 269829 76230 269861
rect 75910 269593 75952 269829
rect 76188 269593 76230 269829
rect 75910 269509 76230 269593
rect 75910 269273 75952 269509
rect 76188 269273 76230 269509
rect 75910 269241 76230 269273
rect 81840 269829 82160 269861
rect 81840 269593 81882 269829
rect 82118 269593 82160 269829
rect 81840 269509 82160 269593
rect 81840 269273 81882 269509
rect 82118 269273 82160 269509
rect 81840 269241 82160 269273
rect 87771 269829 88091 269861
rect 87771 269593 87813 269829
rect 88049 269593 88091 269829
rect 87771 269509 88091 269593
rect 87771 269273 87813 269509
rect 88049 269273 88091 269509
rect 87771 269241 88091 269273
rect 103910 269829 104230 269861
rect 103910 269593 103952 269829
rect 104188 269593 104230 269829
rect 103910 269509 104230 269593
rect 103910 269273 103952 269509
rect 104188 269273 104230 269509
rect 103910 269241 104230 269273
rect 109840 269829 110160 269861
rect 109840 269593 109882 269829
rect 110118 269593 110160 269829
rect 109840 269509 110160 269593
rect 109840 269273 109882 269509
rect 110118 269273 110160 269509
rect 109840 269241 110160 269273
rect 115771 269829 116091 269861
rect 115771 269593 115813 269829
rect 116049 269593 116091 269829
rect 115771 269509 116091 269593
rect 115771 269273 115813 269509
rect 116049 269273 116091 269509
rect 115771 269241 116091 269273
rect 131910 269829 132230 269861
rect 131910 269593 131952 269829
rect 132188 269593 132230 269829
rect 131910 269509 132230 269593
rect 131910 269273 131952 269509
rect 132188 269273 132230 269509
rect 131910 269241 132230 269273
rect 137840 269829 138160 269861
rect 137840 269593 137882 269829
rect 138118 269593 138160 269829
rect 137840 269509 138160 269593
rect 137840 269273 137882 269509
rect 138118 269273 138160 269509
rect 137840 269241 138160 269273
rect 143771 269829 144091 269861
rect 143771 269593 143813 269829
rect 144049 269593 144091 269829
rect 143771 269509 144091 269593
rect 143771 269273 143813 269509
rect 144049 269273 144091 269509
rect 143771 269241 144091 269273
rect 159910 269829 160230 269861
rect 159910 269593 159952 269829
rect 160188 269593 160230 269829
rect 159910 269509 160230 269593
rect 159910 269273 159952 269509
rect 160188 269273 160230 269509
rect 159910 269241 160230 269273
rect 165840 269829 166160 269861
rect 165840 269593 165882 269829
rect 166118 269593 166160 269829
rect 165840 269509 166160 269593
rect 165840 269273 165882 269509
rect 166118 269273 166160 269509
rect 165840 269241 166160 269273
rect 171771 269829 172091 269861
rect 171771 269593 171813 269829
rect 172049 269593 172091 269829
rect 171771 269509 172091 269593
rect 171771 269273 171813 269509
rect 172049 269273 172091 269509
rect 171771 269241 172091 269273
rect 187910 269829 188230 269861
rect 187910 269593 187952 269829
rect 188188 269593 188230 269829
rect 187910 269509 188230 269593
rect 187910 269273 187952 269509
rect 188188 269273 188230 269509
rect 187910 269241 188230 269273
rect 193840 269829 194160 269861
rect 193840 269593 193882 269829
rect 194118 269593 194160 269829
rect 193840 269509 194160 269593
rect 193840 269273 193882 269509
rect 194118 269273 194160 269509
rect 193840 269241 194160 269273
rect 199771 269829 200091 269861
rect 199771 269593 199813 269829
rect 200049 269593 200091 269829
rect 199771 269509 200091 269593
rect 199771 269273 199813 269509
rect 200049 269273 200091 269509
rect 199771 269241 200091 269273
rect 215910 269829 216230 269861
rect 215910 269593 215952 269829
rect 216188 269593 216230 269829
rect 215910 269509 216230 269593
rect 215910 269273 215952 269509
rect 216188 269273 216230 269509
rect 215910 269241 216230 269273
rect 221840 269829 222160 269861
rect 221840 269593 221882 269829
rect 222118 269593 222160 269829
rect 221840 269509 222160 269593
rect 221840 269273 221882 269509
rect 222118 269273 222160 269509
rect 221840 269241 222160 269273
rect 227771 269829 228091 269861
rect 227771 269593 227813 269829
rect 228049 269593 228091 269829
rect 227771 269509 228091 269593
rect 227771 269273 227813 269509
rect 228049 269273 228091 269509
rect 227771 269241 228091 269273
rect 243910 269829 244230 269861
rect 243910 269593 243952 269829
rect 244188 269593 244230 269829
rect 243910 269509 244230 269593
rect 243910 269273 243952 269509
rect 244188 269273 244230 269509
rect 243910 269241 244230 269273
rect 249840 269829 250160 269861
rect 249840 269593 249882 269829
rect 250118 269593 250160 269829
rect 249840 269509 250160 269593
rect 249840 269273 249882 269509
rect 250118 269273 250160 269509
rect 249840 269241 250160 269273
rect 255771 269829 256091 269861
rect 255771 269593 255813 269829
rect 256049 269593 256091 269829
rect 255771 269509 256091 269593
rect 255771 269273 255813 269509
rect 256049 269273 256091 269509
rect 255771 269241 256091 269273
rect 271910 269829 272230 269861
rect 271910 269593 271952 269829
rect 272188 269593 272230 269829
rect 271910 269509 272230 269593
rect 271910 269273 271952 269509
rect 272188 269273 272230 269509
rect 271910 269241 272230 269273
rect 277840 269829 278160 269861
rect 277840 269593 277882 269829
rect 278118 269593 278160 269829
rect 277840 269509 278160 269593
rect 277840 269273 277882 269509
rect 278118 269273 278160 269509
rect 277840 269241 278160 269273
rect 283771 269829 284091 269861
rect 283771 269593 283813 269829
rect 284049 269593 284091 269829
rect 283771 269509 284091 269593
rect 283771 269273 283813 269509
rect 284049 269273 284091 269509
rect 283771 269241 284091 269273
rect 299910 269829 300230 269861
rect 299910 269593 299952 269829
rect 300188 269593 300230 269829
rect 299910 269509 300230 269593
rect 299910 269273 299952 269509
rect 300188 269273 300230 269509
rect 299910 269241 300230 269273
rect 305840 269829 306160 269861
rect 305840 269593 305882 269829
rect 306118 269593 306160 269829
rect 305840 269509 306160 269593
rect 305840 269273 305882 269509
rect 306118 269273 306160 269509
rect 305840 269241 306160 269273
rect 311771 269829 312091 269861
rect 311771 269593 311813 269829
rect 312049 269593 312091 269829
rect 311771 269509 312091 269593
rect 311771 269273 311813 269509
rect 312049 269273 312091 269509
rect 311771 269241 312091 269273
rect 327910 269829 328230 269861
rect 327910 269593 327952 269829
rect 328188 269593 328230 269829
rect 327910 269509 328230 269593
rect 327910 269273 327952 269509
rect 328188 269273 328230 269509
rect 327910 269241 328230 269273
rect 333840 269829 334160 269861
rect 333840 269593 333882 269829
rect 334118 269593 334160 269829
rect 333840 269509 334160 269593
rect 333840 269273 333882 269509
rect 334118 269273 334160 269509
rect 333840 269241 334160 269273
rect 339771 269829 340091 269861
rect 339771 269593 339813 269829
rect 340049 269593 340091 269829
rect 339771 269509 340091 269593
rect 339771 269273 339813 269509
rect 340049 269273 340091 269509
rect 339771 269241 340091 269273
rect 355910 269829 356230 269861
rect 355910 269593 355952 269829
rect 356188 269593 356230 269829
rect 355910 269509 356230 269593
rect 355910 269273 355952 269509
rect 356188 269273 356230 269509
rect 355910 269241 356230 269273
rect 361840 269829 362160 269861
rect 361840 269593 361882 269829
rect 362118 269593 362160 269829
rect 361840 269509 362160 269593
rect 361840 269273 361882 269509
rect 362118 269273 362160 269509
rect 361840 269241 362160 269273
rect 367771 269829 368091 269861
rect 367771 269593 367813 269829
rect 368049 269593 368091 269829
rect 367771 269509 368091 269593
rect 367771 269273 367813 269509
rect 368049 269273 368091 269509
rect 367771 269241 368091 269273
rect 383910 269829 384230 269861
rect 383910 269593 383952 269829
rect 384188 269593 384230 269829
rect 383910 269509 384230 269593
rect 383910 269273 383952 269509
rect 384188 269273 384230 269509
rect 383910 269241 384230 269273
rect 389840 269829 390160 269861
rect 389840 269593 389882 269829
rect 390118 269593 390160 269829
rect 389840 269509 390160 269593
rect 389840 269273 389882 269509
rect 390118 269273 390160 269509
rect 389840 269241 390160 269273
rect 395771 269829 396091 269861
rect 395771 269593 395813 269829
rect 396049 269593 396091 269829
rect 395771 269509 396091 269593
rect 395771 269273 395813 269509
rect 396049 269273 396091 269509
rect 395771 269241 396091 269273
rect 411910 269829 412230 269861
rect 411910 269593 411952 269829
rect 412188 269593 412230 269829
rect 411910 269509 412230 269593
rect 411910 269273 411952 269509
rect 412188 269273 412230 269509
rect 411910 269241 412230 269273
rect 417840 269829 418160 269861
rect 417840 269593 417882 269829
rect 418118 269593 418160 269829
rect 417840 269509 418160 269593
rect 417840 269273 417882 269509
rect 418118 269273 418160 269509
rect 417840 269241 418160 269273
rect 423771 269829 424091 269861
rect 423771 269593 423813 269829
rect 424049 269593 424091 269829
rect 423771 269509 424091 269593
rect 423771 269273 423813 269509
rect 424049 269273 424091 269509
rect 423771 269241 424091 269273
rect 439910 269829 440230 269861
rect 439910 269593 439952 269829
rect 440188 269593 440230 269829
rect 439910 269509 440230 269593
rect 439910 269273 439952 269509
rect 440188 269273 440230 269509
rect 439910 269241 440230 269273
rect 445840 269829 446160 269861
rect 445840 269593 445882 269829
rect 446118 269593 446160 269829
rect 445840 269509 446160 269593
rect 445840 269273 445882 269509
rect 446118 269273 446160 269509
rect 445840 269241 446160 269273
rect 451771 269829 452091 269861
rect 451771 269593 451813 269829
rect 452049 269593 452091 269829
rect 451771 269509 452091 269593
rect 451771 269273 451813 269509
rect 452049 269273 452091 269509
rect 451771 269241 452091 269273
rect 467910 269829 468230 269861
rect 467910 269593 467952 269829
rect 468188 269593 468230 269829
rect 467910 269509 468230 269593
rect 467910 269273 467952 269509
rect 468188 269273 468230 269509
rect 467910 269241 468230 269273
rect 473840 269829 474160 269861
rect 473840 269593 473882 269829
rect 474118 269593 474160 269829
rect 473840 269509 474160 269593
rect 473840 269273 473882 269509
rect 474118 269273 474160 269509
rect 473840 269241 474160 269273
rect 479771 269829 480091 269861
rect 479771 269593 479813 269829
rect 480049 269593 480091 269829
rect 479771 269509 480091 269593
rect 479771 269273 479813 269509
rect 480049 269273 480091 269509
rect 479771 269241 480091 269273
rect 495910 269829 496230 269861
rect 495910 269593 495952 269829
rect 496188 269593 496230 269829
rect 495910 269509 496230 269593
rect 495910 269273 495952 269509
rect 496188 269273 496230 269509
rect 495910 269241 496230 269273
rect 501840 269829 502160 269861
rect 501840 269593 501882 269829
rect 502118 269593 502160 269829
rect 501840 269509 502160 269593
rect 501840 269273 501882 269509
rect 502118 269273 502160 269509
rect 501840 269241 502160 269273
rect 507771 269829 508091 269861
rect 507771 269593 507813 269829
rect 508049 269593 508091 269829
rect 507771 269509 508091 269593
rect 507771 269273 507813 269509
rect 508049 269273 508091 269509
rect 507771 269241 508091 269273
rect 523910 269829 524230 269861
rect 523910 269593 523952 269829
rect 524188 269593 524230 269829
rect 523910 269509 524230 269593
rect 523910 269273 523952 269509
rect 524188 269273 524230 269509
rect 523910 269241 524230 269273
rect 529840 269829 530160 269861
rect 529840 269593 529882 269829
rect 530118 269593 530160 269829
rect 529840 269509 530160 269593
rect 529840 269273 529882 269509
rect 530118 269273 530160 269509
rect 529840 269241 530160 269273
rect 535771 269829 536091 269861
rect 535771 269593 535813 269829
rect 536049 269593 536091 269829
rect 535771 269509 536091 269593
rect 535771 269273 535813 269509
rect 536049 269273 536091 269509
rect 535771 269241 536091 269273
rect 551910 269829 552230 269861
rect 551910 269593 551952 269829
rect 552188 269593 552230 269829
rect 551910 269509 552230 269593
rect 551910 269273 551952 269509
rect 552188 269273 552230 269509
rect 551910 269241 552230 269273
rect 557840 269829 558160 269861
rect 557840 269593 557882 269829
rect 558118 269593 558160 269829
rect 557840 269509 558160 269593
rect 557840 269273 557882 269509
rect 558118 269273 558160 269509
rect 557840 269241 558160 269273
rect 563771 269829 564091 269861
rect 563771 269593 563813 269829
rect 564049 269593 564091 269829
rect 563771 269509 564091 269593
rect 563771 269273 563813 269509
rect 564049 269273 564091 269509
rect 563771 269241 564091 269273
rect 573494 269829 574114 296273
rect 573494 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 574114 269829
rect 573494 269509 574114 269593
rect 573494 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 574114 269509
rect 22874 266454 23194 266486
rect 22874 266218 22916 266454
rect 23152 266218 23194 266454
rect 22874 266134 23194 266218
rect 22874 265898 22916 266134
rect 23152 265898 23194 266134
rect 22874 265866 23194 265898
rect 28805 266454 29125 266486
rect 28805 266218 28847 266454
rect 29083 266218 29125 266454
rect 28805 266134 29125 266218
rect 28805 265898 28847 266134
rect 29083 265898 29125 266134
rect 28805 265866 29125 265898
rect 50874 266454 51194 266486
rect 50874 266218 50916 266454
rect 51152 266218 51194 266454
rect 50874 266134 51194 266218
rect 50874 265898 50916 266134
rect 51152 265898 51194 266134
rect 50874 265866 51194 265898
rect 56805 266454 57125 266486
rect 56805 266218 56847 266454
rect 57083 266218 57125 266454
rect 56805 266134 57125 266218
rect 56805 265898 56847 266134
rect 57083 265898 57125 266134
rect 56805 265866 57125 265898
rect 78874 266454 79194 266486
rect 78874 266218 78916 266454
rect 79152 266218 79194 266454
rect 78874 266134 79194 266218
rect 78874 265898 78916 266134
rect 79152 265898 79194 266134
rect 78874 265866 79194 265898
rect 84805 266454 85125 266486
rect 84805 266218 84847 266454
rect 85083 266218 85125 266454
rect 84805 266134 85125 266218
rect 84805 265898 84847 266134
rect 85083 265898 85125 266134
rect 84805 265866 85125 265898
rect 106874 266454 107194 266486
rect 106874 266218 106916 266454
rect 107152 266218 107194 266454
rect 106874 266134 107194 266218
rect 106874 265898 106916 266134
rect 107152 265898 107194 266134
rect 106874 265866 107194 265898
rect 112805 266454 113125 266486
rect 112805 266218 112847 266454
rect 113083 266218 113125 266454
rect 112805 266134 113125 266218
rect 112805 265898 112847 266134
rect 113083 265898 113125 266134
rect 112805 265866 113125 265898
rect 134874 266454 135194 266486
rect 134874 266218 134916 266454
rect 135152 266218 135194 266454
rect 134874 266134 135194 266218
rect 134874 265898 134916 266134
rect 135152 265898 135194 266134
rect 134874 265866 135194 265898
rect 140805 266454 141125 266486
rect 140805 266218 140847 266454
rect 141083 266218 141125 266454
rect 140805 266134 141125 266218
rect 140805 265898 140847 266134
rect 141083 265898 141125 266134
rect 140805 265866 141125 265898
rect 162874 266454 163194 266486
rect 162874 266218 162916 266454
rect 163152 266218 163194 266454
rect 162874 266134 163194 266218
rect 162874 265898 162916 266134
rect 163152 265898 163194 266134
rect 162874 265866 163194 265898
rect 168805 266454 169125 266486
rect 168805 266218 168847 266454
rect 169083 266218 169125 266454
rect 168805 266134 169125 266218
rect 168805 265898 168847 266134
rect 169083 265898 169125 266134
rect 168805 265866 169125 265898
rect 190874 266454 191194 266486
rect 190874 266218 190916 266454
rect 191152 266218 191194 266454
rect 190874 266134 191194 266218
rect 190874 265898 190916 266134
rect 191152 265898 191194 266134
rect 190874 265866 191194 265898
rect 196805 266454 197125 266486
rect 196805 266218 196847 266454
rect 197083 266218 197125 266454
rect 196805 266134 197125 266218
rect 196805 265898 196847 266134
rect 197083 265898 197125 266134
rect 196805 265866 197125 265898
rect 218874 266454 219194 266486
rect 218874 266218 218916 266454
rect 219152 266218 219194 266454
rect 218874 266134 219194 266218
rect 218874 265898 218916 266134
rect 219152 265898 219194 266134
rect 218874 265866 219194 265898
rect 224805 266454 225125 266486
rect 224805 266218 224847 266454
rect 225083 266218 225125 266454
rect 224805 266134 225125 266218
rect 224805 265898 224847 266134
rect 225083 265898 225125 266134
rect 224805 265866 225125 265898
rect 246874 266454 247194 266486
rect 246874 266218 246916 266454
rect 247152 266218 247194 266454
rect 246874 266134 247194 266218
rect 246874 265898 246916 266134
rect 247152 265898 247194 266134
rect 246874 265866 247194 265898
rect 252805 266454 253125 266486
rect 252805 266218 252847 266454
rect 253083 266218 253125 266454
rect 252805 266134 253125 266218
rect 252805 265898 252847 266134
rect 253083 265898 253125 266134
rect 252805 265866 253125 265898
rect 274874 266454 275194 266486
rect 274874 266218 274916 266454
rect 275152 266218 275194 266454
rect 274874 266134 275194 266218
rect 274874 265898 274916 266134
rect 275152 265898 275194 266134
rect 274874 265866 275194 265898
rect 280805 266454 281125 266486
rect 280805 266218 280847 266454
rect 281083 266218 281125 266454
rect 280805 266134 281125 266218
rect 280805 265898 280847 266134
rect 281083 265898 281125 266134
rect 280805 265866 281125 265898
rect 302874 266454 303194 266486
rect 302874 266218 302916 266454
rect 303152 266218 303194 266454
rect 302874 266134 303194 266218
rect 302874 265898 302916 266134
rect 303152 265898 303194 266134
rect 302874 265866 303194 265898
rect 308805 266454 309125 266486
rect 308805 266218 308847 266454
rect 309083 266218 309125 266454
rect 308805 266134 309125 266218
rect 308805 265898 308847 266134
rect 309083 265898 309125 266134
rect 308805 265866 309125 265898
rect 330874 266454 331194 266486
rect 330874 266218 330916 266454
rect 331152 266218 331194 266454
rect 330874 266134 331194 266218
rect 330874 265898 330916 266134
rect 331152 265898 331194 266134
rect 330874 265866 331194 265898
rect 336805 266454 337125 266486
rect 336805 266218 336847 266454
rect 337083 266218 337125 266454
rect 336805 266134 337125 266218
rect 336805 265898 336847 266134
rect 337083 265898 337125 266134
rect 336805 265866 337125 265898
rect 358874 266454 359194 266486
rect 358874 266218 358916 266454
rect 359152 266218 359194 266454
rect 358874 266134 359194 266218
rect 358874 265898 358916 266134
rect 359152 265898 359194 266134
rect 358874 265866 359194 265898
rect 364805 266454 365125 266486
rect 364805 266218 364847 266454
rect 365083 266218 365125 266454
rect 364805 266134 365125 266218
rect 364805 265898 364847 266134
rect 365083 265898 365125 266134
rect 364805 265866 365125 265898
rect 386874 266454 387194 266486
rect 386874 266218 386916 266454
rect 387152 266218 387194 266454
rect 386874 266134 387194 266218
rect 386874 265898 386916 266134
rect 387152 265898 387194 266134
rect 386874 265866 387194 265898
rect 392805 266454 393125 266486
rect 392805 266218 392847 266454
rect 393083 266218 393125 266454
rect 392805 266134 393125 266218
rect 392805 265898 392847 266134
rect 393083 265898 393125 266134
rect 392805 265866 393125 265898
rect 414874 266454 415194 266486
rect 414874 266218 414916 266454
rect 415152 266218 415194 266454
rect 414874 266134 415194 266218
rect 414874 265898 414916 266134
rect 415152 265898 415194 266134
rect 414874 265866 415194 265898
rect 420805 266454 421125 266486
rect 420805 266218 420847 266454
rect 421083 266218 421125 266454
rect 420805 266134 421125 266218
rect 420805 265898 420847 266134
rect 421083 265898 421125 266134
rect 420805 265866 421125 265898
rect 442874 266454 443194 266486
rect 442874 266218 442916 266454
rect 443152 266218 443194 266454
rect 442874 266134 443194 266218
rect 442874 265898 442916 266134
rect 443152 265898 443194 266134
rect 442874 265866 443194 265898
rect 448805 266454 449125 266486
rect 448805 266218 448847 266454
rect 449083 266218 449125 266454
rect 448805 266134 449125 266218
rect 448805 265898 448847 266134
rect 449083 265898 449125 266134
rect 448805 265866 449125 265898
rect 470874 266454 471194 266486
rect 470874 266218 470916 266454
rect 471152 266218 471194 266454
rect 470874 266134 471194 266218
rect 470874 265898 470916 266134
rect 471152 265898 471194 266134
rect 470874 265866 471194 265898
rect 476805 266454 477125 266486
rect 476805 266218 476847 266454
rect 477083 266218 477125 266454
rect 476805 266134 477125 266218
rect 476805 265898 476847 266134
rect 477083 265898 477125 266134
rect 476805 265866 477125 265898
rect 498874 266454 499194 266486
rect 498874 266218 498916 266454
rect 499152 266218 499194 266454
rect 498874 266134 499194 266218
rect 498874 265898 498916 266134
rect 499152 265898 499194 266134
rect 498874 265866 499194 265898
rect 504805 266454 505125 266486
rect 504805 266218 504847 266454
rect 505083 266218 505125 266454
rect 504805 266134 505125 266218
rect 504805 265898 504847 266134
rect 505083 265898 505125 266134
rect 504805 265866 505125 265898
rect 526874 266454 527194 266486
rect 526874 266218 526916 266454
rect 527152 266218 527194 266454
rect 526874 266134 527194 266218
rect 526874 265898 526916 266134
rect 527152 265898 527194 266134
rect 526874 265866 527194 265898
rect 532805 266454 533125 266486
rect 532805 266218 532847 266454
rect 533083 266218 533125 266454
rect 532805 266134 533125 266218
rect 532805 265898 532847 266134
rect 533083 265898 533125 266134
rect 532805 265866 533125 265898
rect 554874 266454 555194 266486
rect 554874 266218 554916 266454
rect 555152 266218 555194 266454
rect 554874 266134 555194 266218
rect 554874 265898 554916 266134
rect 555152 265898 555194 266134
rect 554874 265866 555194 265898
rect 560805 266454 561125 266486
rect 560805 266218 560847 266454
rect 561083 266218 561125 266454
rect 560805 266134 561125 266218
rect 560805 265898 560847 266134
rect 561083 265898 561125 266134
rect 560805 265866 561125 265898
rect -2006 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 -1386 242829
rect -2006 242509 -1386 242593
rect -2006 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 -1386 242509
rect -2006 215829 -1386 242273
rect 19910 242829 20230 242861
rect 19910 242593 19952 242829
rect 20188 242593 20230 242829
rect 19910 242509 20230 242593
rect 19910 242273 19952 242509
rect 20188 242273 20230 242509
rect 19910 242241 20230 242273
rect 25840 242829 26160 242861
rect 25840 242593 25882 242829
rect 26118 242593 26160 242829
rect 25840 242509 26160 242593
rect 25840 242273 25882 242509
rect 26118 242273 26160 242509
rect 25840 242241 26160 242273
rect 31771 242829 32091 242861
rect 31771 242593 31813 242829
rect 32049 242593 32091 242829
rect 31771 242509 32091 242593
rect 31771 242273 31813 242509
rect 32049 242273 32091 242509
rect 31771 242241 32091 242273
rect 47910 242829 48230 242861
rect 47910 242593 47952 242829
rect 48188 242593 48230 242829
rect 47910 242509 48230 242593
rect 47910 242273 47952 242509
rect 48188 242273 48230 242509
rect 47910 242241 48230 242273
rect 53840 242829 54160 242861
rect 53840 242593 53882 242829
rect 54118 242593 54160 242829
rect 53840 242509 54160 242593
rect 53840 242273 53882 242509
rect 54118 242273 54160 242509
rect 53840 242241 54160 242273
rect 59771 242829 60091 242861
rect 59771 242593 59813 242829
rect 60049 242593 60091 242829
rect 59771 242509 60091 242593
rect 59771 242273 59813 242509
rect 60049 242273 60091 242509
rect 59771 242241 60091 242273
rect 75910 242829 76230 242861
rect 75910 242593 75952 242829
rect 76188 242593 76230 242829
rect 75910 242509 76230 242593
rect 75910 242273 75952 242509
rect 76188 242273 76230 242509
rect 75910 242241 76230 242273
rect 81840 242829 82160 242861
rect 81840 242593 81882 242829
rect 82118 242593 82160 242829
rect 81840 242509 82160 242593
rect 81840 242273 81882 242509
rect 82118 242273 82160 242509
rect 81840 242241 82160 242273
rect 87771 242829 88091 242861
rect 87771 242593 87813 242829
rect 88049 242593 88091 242829
rect 87771 242509 88091 242593
rect 87771 242273 87813 242509
rect 88049 242273 88091 242509
rect 87771 242241 88091 242273
rect 103910 242829 104230 242861
rect 103910 242593 103952 242829
rect 104188 242593 104230 242829
rect 103910 242509 104230 242593
rect 103910 242273 103952 242509
rect 104188 242273 104230 242509
rect 103910 242241 104230 242273
rect 109840 242829 110160 242861
rect 109840 242593 109882 242829
rect 110118 242593 110160 242829
rect 109840 242509 110160 242593
rect 109840 242273 109882 242509
rect 110118 242273 110160 242509
rect 109840 242241 110160 242273
rect 115771 242829 116091 242861
rect 115771 242593 115813 242829
rect 116049 242593 116091 242829
rect 115771 242509 116091 242593
rect 115771 242273 115813 242509
rect 116049 242273 116091 242509
rect 115771 242241 116091 242273
rect 131910 242829 132230 242861
rect 131910 242593 131952 242829
rect 132188 242593 132230 242829
rect 131910 242509 132230 242593
rect 131910 242273 131952 242509
rect 132188 242273 132230 242509
rect 131910 242241 132230 242273
rect 137840 242829 138160 242861
rect 137840 242593 137882 242829
rect 138118 242593 138160 242829
rect 137840 242509 138160 242593
rect 137840 242273 137882 242509
rect 138118 242273 138160 242509
rect 137840 242241 138160 242273
rect 143771 242829 144091 242861
rect 143771 242593 143813 242829
rect 144049 242593 144091 242829
rect 143771 242509 144091 242593
rect 143771 242273 143813 242509
rect 144049 242273 144091 242509
rect 143771 242241 144091 242273
rect 159910 242829 160230 242861
rect 159910 242593 159952 242829
rect 160188 242593 160230 242829
rect 159910 242509 160230 242593
rect 159910 242273 159952 242509
rect 160188 242273 160230 242509
rect 159910 242241 160230 242273
rect 165840 242829 166160 242861
rect 165840 242593 165882 242829
rect 166118 242593 166160 242829
rect 165840 242509 166160 242593
rect 165840 242273 165882 242509
rect 166118 242273 166160 242509
rect 165840 242241 166160 242273
rect 171771 242829 172091 242861
rect 171771 242593 171813 242829
rect 172049 242593 172091 242829
rect 171771 242509 172091 242593
rect 171771 242273 171813 242509
rect 172049 242273 172091 242509
rect 171771 242241 172091 242273
rect 187910 242829 188230 242861
rect 187910 242593 187952 242829
rect 188188 242593 188230 242829
rect 187910 242509 188230 242593
rect 187910 242273 187952 242509
rect 188188 242273 188230 242509
rect 187910 242241 188230 242273
rect 193840 242829 194160 242861
rect 193840 242593 193882 242829
rect 194118 242593 194160 242829
rect 193840 242509 194160 242593
rect 193840 242273 193882 242509
rect 194118 242273 194160 242509
rect 193840 242241 194160 242273
rect 199771 242829 200091 242861
rect 199771 242593 199813 242829
rect 200049 242593 200091 242829
rect 199771 242509 200091 242593
rect 199771 242273 199813 242509
rect 200049 242273 200091 242509
rect 199771 242241 200091 242273
rect 215910 242829 216230 242861
rect 215910 242593 215952 242829
rect 216188 242593 216230 242829
rect 215910 242509 216230 242593
rect 215910 242273 215952 242509
rect 216188 242273 216230 242509
rect 215910 242241 216230 242273
rect 221840 242829 222160 242861
rect 221840 242593 221882 242829
rect 222118 242593 222160 242829
rect 221840 242509 222160 242593
rect 221840 242273 221882 242509
rect 222118 242273 222160 242509
rect 221840 242241 222160 242273
rect 227771 242829 228091 242861
rect 227771 242593 227813 242829
rect 228049 242593 228091 242829
rect 227771 242509 228091 242593
rect 227771 242273 227813 242509
rect 228049 242273 228091 242509
rect 227771 242241 228091 242273
rect 243910 242829 244230 242861
rect 243910 242593 243952 242829
rect 244188 242593 244230 242829
rect 243910 242509 244230 242593
rect 243910 242273 243952 242509
rect 244188 242273 244230 242509
rect 243910 242241 244230 242273
rect 249840 242829 250160 242861
rect 249840 242593 249882 242829
rect 250118 242593 250160 242829
rect 249840 242509 250160 242593
rect 249840 242273 249882 242509
rect 250118 242273 250160 242509
rect 249840 242241 250160 242273
rect 255771 242829 256091 242861
rect 255771 242593 255813 242829
rect 256049 242593 256091 242829
rect 255771 242509 256091 242593
rect 255771 242273 255813 242509
rect 256049 242273 256091 242509
rect 255771 242241 256091 242273
rect 271910 242829 272230 242861
rect 271910 242593 271952 242829
rect 272188 242593 272230 242829
rect 271910 242509 272230 242593
rect 271910 242273 271952 242509
rect 272188 242273 272230 242509
rect 271910 242241 272230 242273
rect 277840 242829 278160 242861
rect 277840 242593 277882 242829
rect 278118 242593 278160 242829
rect 277840 242509 278160 242593
rect 277840 242273 277882 242509
rect 278118 242273 278160 242509
rect 277840 242241 278160 242273
rect 283771 242829 284091 242861
rect 283771 242593 283813 242829
rect 284049 242593 284091 242829
rect 283771 242509 284091 242593
rect 283771 242273 283813 242509
rect 284049 242273 284091 242509
rect 283771 242241 284091 242273
rect 299910 242829 300230 242861
rect 299910 242593 299952 242829
rect 300188 242593 300230 242829
rect 299910 242509 300230 242593
rect 299910 242273 299952 242509
rect 300188 242273 300230 242509
rect 299910 242241 300230 242273
rect 305840 242829 306160 242861
rect 305840 242593 305882 242829
rect 306118 242593 306160 242829
rect 305840 242509 306160 242593
rect 305840 242273 305882 242509
rect 306118 242273 306160 242509
rect 305840 242241 306160 242273
rect 311771 242829 312091 242861
rect 311771 242593 311813 242829
rect 312049 242593 312091 242829
rect 311771 242509 312091 242593
rect 311771 242273 311813 242509
rect 312049 242273 312091 242509
rect 311771 242241 312091 242273
rect 327910 242829 328230 242861
rect 327910 242593 327952 242829
rect 328188 242593 328230 242829
rect 327910 242509 328230 242593
rect 327910 242273 327952 242509
rect 328188 242273 328230 242509
rect 327910 242241 328230 242273
rect 333840 242829 334160 242861
rect 333840 242593 333882 242829
rect 334118 242593 334160 242829
rect 333840 242509 334160 242593
rect 333840 242273 333882 242509
rect 334118 242273 334160 242509
rect 333840 242241 334160 242273
rect 339771 242829 340091 242861
rect 339771 242593 339813 242829
rect 340049 242593 340091 242829
rect 339771 242509 340091 242593
rect 339771 242273 339813 242509
rect 340049 242273 340091 242509
rect 339771 242241 340091 242273
rect 355910 242829 356230 242861
rect 355910 242593 355952 242829
rect 356188 242593 356230 242829
rect 355910 242509 356230 242593
rect 355910 242273 355952 242509
rect 356188 242273 356230 242509
rect 355910 242241 356230 242273
rect 361840 242829 362160 242861
rect 361840 242593 361882 242829
rect 362118 242593 362160 242829
rect 361840 242509 362160 242593
rect 361840 242273 361882 242509
rect 362118 242273 362160 242509
rect 361840 242241 362160 242273
rect 367771 242829 368091 242861
rect 367771 242593 367813 242829
rect 368049 242593 368091 242829
rect 367771 242509 368091 242593
rect 367771 242273 367813 242509
rect 368049 242273 368091 242509
rect 367771 242241 368091 242273
rect 383910 242829 384230 242861
rect 383910 242593 383952 242829
rect 384188 242593 384230 242829
rect 383910 242509 384230 242593
rect 383910 242273 383952 242509
rect 384188 242273 384230 242509
rect 383910 242241 384230 242273
rect 389840 242829 390160 242861
rect 389840 242593 389882 242829
rect 390118 242593 390160 242829
rect 389840 242509 390160 242593
rect 389840 242273 389882 242509
rect 390118 242273 390160 242509
rect 389840 242241 390160 242273
rect 395771 242829 396091 242861
rect 395771 242593 395813 242829
rect 396049 242593 396091 242829
rect 395771 242509 396091 242593
rect 395771 242273 395813 242509
rect 396049 242273 396091 242509
rect 395771 242241 396091 242273
rect 411910 242829 412230 242861
rect 411910 242593 411952 242829
rect 412188 242593 412230 242829
rect 411910 242509 412230 242593
rect 411910 242273 411952 242509
rect 412188 242273 412230 242509
rect 411910 242241 412230 242273
rect 417840 242829 418160 242861
rect 417840 242593 417882 242829
rect 418118 242593 418160 242829
rect 417840 242509 418160 242593
rect 417840 242273 417882 242509
rect 418118 242273 418160 242509
rect 417840 242241 418160 242273
rect 423771 242829 424091 242861
rect 423771 242593 423813 242829
rect 424049 242593 424091 242829
rect 423771 242509 424091 242593
rect 423771 242273 423813 242509
rect 424049 242273 424091 242509
rect 423771 242241 424091 242273
rect 439910 242829 440230 242861
rect 439910 242593 439952 242829
rect 440188 242593 440230 242829
rect 439910 242509 440230 242593
rect 439910 242273 439952 242509
rect 440188 242273 440230 242509
rect 439910 242241 440230 242273
rect 445840 242829 446160 242861
rect 445840 242593 445882 242829
rect 446118 242593 446160 242829
rect 445840 242509 446160 242593
rect 445840 242273 445882 242509
rect 446118 242273 446160 242509
rect 445840 242241 446160 242273
rect 451771 242829 452091 242861
rect 451771 242593 451813 242829
rect 452049 242593 452091 242829
rect 451771 242509 452091 242593
rect 451771 242273 451813 242509
rect 452049 242273 452091 242509
rect 451771 242241 452091 242273
rect 467910 242829 468230 242861
rect 467910 242593 467952 242829
rect 468188 242593 468230 242829
rect 467910 242509 468230 242593
rect 467910 242273 467952 242509
rect 468188 242273 468230 242509
rect 467910 242241 468230 242273
rect 473840 242829 474160 242861
rect 473840 242593 473882 242829
rect 474118 242593 474160 242829
rect 473840 242509 474160 242593
rect 473840 242273 473882 242509
rect 474118 242273 474160 242509
rect 473840 242241 474160 242273
rect 479771 242829 480091 242861
rect 479771 242593 479813 242829
rect 480049 242593 480091 242829
rect 479771 242509 480091 242593
rect 479771 242273 479813 242509
rect 480049 242273 480091 242509
rect 479771 242241 480091 242273
rect 495910 242829 496230 242861
rect 495910 242593 495952 242829
rect 496188 242593 496230 242829
rect 495910 242509 496230 242593
rect 495910 242273 495952 242509
rect 496188 242273 496230 242509
rect 495910 242241 496230 242273
rect 501840 242829 502160 242861
rect 501840 242593 501882 242829
rect 502118 242593 502160 242829
rect 501840 242509 502160 242593
rect 501840 242273 501882 242509
rect 502118 242273 502160 242509
rect 501840 242241 502160 242273
rect 507771 242829 508091 242861
rect 507771 242593 507813 242829
rect 508049 242593 508091 242829
rect 507771 242509 508091 242593
rect 507771 242273 507813 242509
rect 508049 242273 508091 242509
rect 507771 242241 508091 242273
rect 523910 242829 524230 242861
rect 523910 242593 523952 242829
rect 524188 242593 524230 242829
rect 523910 242509 524230 242593
rect 523910 242273 523952 242509
rect 524188 242273 524230 242509
rect 523910 242241 524230 242273
rect 529840 242829 530160 242861
rect 529840 242593 529882 242829
rect 530118 242593 530160 242829
rect 529840 242509 530160 242593
rect 529840 242273 529882 242509
rect 530118 242273 530160 242509
rect 529840 242241 530160 242273
rect 535771 242829 536091 242861
rect 535771 242593 535813 242829
rect 536049 242593 536091 242829
rect 535771 242509 536091 242593
rect 535771 242273 535813 242509
rect 536049 242273 536091 242509
rect 535771 242241 536091 242273
rect 551910 242829 552230 242861
rect 551910 242593 551952 242829
rect 552188 242593 552230 242829
rect 551910 242509 552230 242593
rect 551910 242273 551952 242509
rect 552188 242273 552230 242509
rect 551910 242241 552230 242273
rect 557840 242829 558160 242861
rect 557840 242593 557882 242829
rect 558118 242593 558160 242829
rect 557840 242509 558160 242593
rect 557840 242273 557882 242509
rect 558118 242273 558160 242509
rect 557840 242241 558160 242273
rect 563771 242829 564091 242861
rect 563771 242593 563813 242829
rect 564049 242593 564091 242829
rect 563771 242509 564091 242593
rect 563771 242273 563813 242509
rect 564049 242273 564091 242509
rect 563771 242241 564091 242273
rect 573494 242829 574114 269273
rect 573494 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 574114 242829
rect 573494 242509 574114 242593
rect 573494 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 574114 242509
rect 22874 239454 23194 239486
rect 22874 239218 22916 239454
rect 23152 239218 23194 239454
rect 22874 239134 23194 239218
rect 22874 238898 22916 239134
rect 23152 238898 23194 239134
rect 22874 238866 23194 238898
rect 28805 239454 29125 239486
rect 28805 239218 28847 239454
rect 29083 239218 29125 239454
rect 28805 239134 29125 239218
rect 28805 238898 28847 239134
rect 29083 238898 29125 239134
rect 28805 238866 29125 238898
rect 50874 239454 51194 239486
rect 50874 239218 50916 239454
rect 51152 239218 51194 239454
rect 50874 239134 51194 239218
rect 50874 238898 50916 239134
rect 51152 238898 51194 239134
rect 50874 238866 51194 238898
rect 56805 239454 57125 239486
rect 56805 239218 56847 239454
rect 57083 239218 57125 239454
rect 56805 239134 57125 239218
rect 56805 238898 56847 239134
rect 57083 238898 57125 239134
rect 56805 238866 57125 238898
rect 78874 239454 79194 239486
rect 78874 239218 78916 239454
rect 79152 239218 79194 239454
rect 78874 239134 79194 239218
rect 78874 238898 78916 239134
rect 79152 238898 79194 239134
rect 78874 238866 79194 238898
rect 84805 239454 85125 239486
rect 84805 239218 84847 239454
rect 85083 239218 85125 239454
rect 84805 239134 85125 239218
rect 84805 238898 84847 239134
rect 85083 238898 85125 239134
rect 84805 238866 85125 238898
rect 106874 239454 107194 239486
rect 106874 239218 106916 239454
rect 107152 239218 107194 239454
rect 106874 239134 107194 239218
rect 106874 238898 106916 239134
rect 107152 238898 107194 239134
rect 106874 238866 107194 238898
rect 112805 239454 113125 239486
rect 112805 239218 112847 239454
rect 113083 239218 113125 239454
rect 112805 239134 113125 239218
rect 112805 238898 112847 239134
rect 113083 238898 113125 239134
rect 112805 238866 113125 238898
rect 134874 239454 135194 239486
rect 134874 239218 134916 239454
rect 135152 239218 135194 239454
rect 134874 239134 135194 239218
rect 134874 238898 134916 239134
rect 135152 238898 135194 239134
rect 134874 238866 135194 238898
rect 140805 239454 141125 239486
rect 140805 239218 140847 239454
rect 141083 239218 141125 239454
rect 140805 239134 141125 239218
rect 140805 238898 140847 239134
rect 141083 238898 141125 239134
rect 140805 238866 141125 238898
rect 162874 239454 163194 239486
rect 162874 239218 162916 239454
rect 163152 239218 163194 239454
rect 162874 239134 163194 239218
rect 162874 238898 162916 239134
rect 163152 238898 163194 239134
rect 162874 238866 163194 238898
rect 168805 239454 169125 239486
rect 168805 239218 168847 239454
rect 169083 239218 169125 239454
rect 168805 239134 169125 239218
rect 168805 238898 168847 239134
rect 169083 238898 169125 239134
rect 168805 238866 169125 238898
rect 190874 239454 191194 239486
rect 190874 239218 190916 239454
rect 191152 239218 191194 239454
rect 190874 239134 191194 239218
rect 190874 238898 190916 239134
rect 191152 238898 191194 239134
rect 190874 238866 191194 238898
rect 196805 239454 197125 239486
rect 196805 239218 196847 239454
rect 197083 239218 197125 239454
rect 196805 239134 197125 239218
rect 196805 238898 196847 239134
rect 197083 238898 197125 239134
rect 196805 238866 197125 238898
rect 218874 239454 219194 239486
rect 218874 239218 218916 239454
rect 219152 239218 219194 239454
rect 218874 239134 219194 239218
rect 218874 238898 218916 239134
rect 219152 238898 219194 239134
rect 218874 238866 219194 238898
rect 224805 239454 225125 239486
rect 224805 239218 224847 239454
rect 225083 239218 225125 239454
rect 224805 239134 225125 239218
rect 224805 238898 224847 239134
rect 225083 238898 225125 239134
rect 224805 238866 225125 238898
rect 246874 239454 247194 239486
rect 246874 239218 246916 239454
rect 247152 239218 247194 239454
rect 246874 239134 247194 239218
rect 246874 238898 246916 239134
rect 247152 238898 247194 239134
rect 246874 238866 247194 238898
rect 252805 239454 253125 239486
rect 252805 239218 252847 239454
rect 253083 239218 253125 239454
rect 252805 239134 253125 239218
rect 252805 238898 252847 239134
rect 253083 238898 253125 239134
rect 252805 238866 253125 238898
rect 274874 239454 275194 239486
rect 274874 239218 274916 239454
rect 275152 239218 275194 239454
rect 274874 239134 275194 239218
rect 274874 238898 274916 239134
rect 275152 238898 275194 239134
rect 274874 238866 275194 238898
rect 280805 239454 281125 239486
rect 280805 239218 280847 239454
rect 281083 239218 281125 239454
rect 280805 239134 281125 239218
rect 280805 238898 280847 239134
rect 281083 238898 281125 239134
rect 280805 238866 281125 238898
rect 302874 239454 303194 239486
rect 302874 239218 302916 239454
rect 303152 239218 303194 239454
rect 302874 239134 303194 239218
rect 302874 238898 302916 239134
rect 303152 238898 303194 239134
rect 302874 238866 303194 238898
rect 308805 239454 309125 239486
rect 308805 239218 308847 239454
rect 309083 239218 309125 239454
rect 308805 239134 309125 239218
rect 308805 238898 308847 239134
rect 309083 238898 309125 239134
rect 308805 238866 309125 238898
rect 330874 239454 331194 239486
rect 330874 239218 330916 239454
rect 331152 239218 331194 239454
rect 330874 239134 331194 239218
rect 330874 238898 330916 239134
rect 331152 238898 331194 239134
rect 330874 238866 331194 238898
rect 336805 239454 337125 239486
rect 336805 239218 336847 239454
rect 337083 239218 337125 239454
rect 336805 239134 337125 239218
rect 336805 238898 336847 239134
rect 337083 238898 337125 239134
rect 336805 238866 337125 238898
rect 358874 239454 359194 239486
rect 358874 239218 358916 239454
rect 359152 239218 359194 239454
rect 358874 239134 359194 239218
rect 358874 238898 358916 239134
rect 359152 238898 359194 239134
rect 358874 238866 359194 238898
rect 364805 239454 365125 239486
rect 364805 239218 364847 239454
rect 365083 239218 365125 239454
rect 364805 239134 365125 239218
rect 364805 238898 364847 239134
rect 365083 238898 365125 239134
rect 364805 238866 365125 238898
rect 386874 239454 387194 239486
rect 386874 239218 386916 239454
rect 387152 239218 387194 239454
rect 386874 239134 387194 239218
rect 386874 238898 386916 239134
rect 387152 238898 387194 239134
rect 386874 238866 387194 238898
rect 392805 239454 393125 239486
rect 392805 239218 392847 239454
rect 393083 239218 393125 239454
rect 392805 239134 393125 239218
rect 392805 238898 392847 239134
rect 393083 238898 393125 239134
rect 392805 238866 393125 238898
rect 414874 239454 415194 239486
rect 414874 239218 414916 239454
rect 415152 239218 415194 239454
rect 414874 239134 415194 239218
rect 414874 238898 414916 239134
rect 415152 238898 415194 239134
rect 414874 238866 415194 238898
rect 420805 239454 421125 239486
rect 420805 239218 420847 239454
rect 421083 239218 421125 239454
rect 420805 239134 421125 239218
rect 420805 238898 420847 239134
rect 421083 238898 421125 239134
rect 420805 238866 421125 238898
rect 442874 239454 443194 239486
rect 442874 239218 442916 239454
rect 443152 239218 443194 239454
rect 442874 239134 443194 239218
rect 442874 238898 442916 239134
rect 443152 238898 443194 239134
rect 442874 238866 443194 238898
rect 448805 239454 449125 239486
rect 448805 239218 448847 239454
rect 449083 239218 449125 239454
rect 448805 239134 449125 239218
rect 448805 238898 448847 239134
rect 449083 238898 449125 239134
rect 448805 238866 449125 238898
rect 470874 239454 471194 239486
rect 470874 239218 470916 239454
rect 471152 239218 471194 239454
rect 470874 239134 471194 239218
rect 470874 238898 470916 239134
rect 471152 238898 471194 239134
rect 470874 238866 471194 238898
rect 476805 239454 477125 239486
rect 476805 239218 476847 239454
rect 477083 239218 477125 239454
rect 476805 239134 477125 239218
rect 476805 238898 476847 239134
rect 477083 238898 477125 239134
rect 476805 238866 477125 238898
rect 498874 239454 499194 239486
rect 498874 239218 498916 239454
rect 499152 239218 499194 239454
rect 498874 239134 499194 239218
rect 498874 238898 498916 239134
rect 499152 238898 499194 239134
rect 498874 238866 499194 238898
rect 504805 239454 505125 239486
rect 504805 239218 504847 239454
rect 505083 239218 505125 239454
rect 504805 239134 505125 239218
rect 504805 238898 504847 239134
rect 505083 238898 505125 239134
rect 504805 238866 505125 238898
rect 526874 239454 527194 239486
rect 526874 239218 526916 239454
rect 527152 239218 527194 239454
rect 526874 239134 527194 239218
rect 526874 238898 526916 239134
rect 527152 238898 527194 239134
rect 526874 238866 527194 238898
rect 532805 239454 533125 239486
rect 532805 239218 532847 239454
rect 533083 239218 533125 239454
rect 532805 239134 533125 239218
rect 532805 238898 532847 239134
rect 533083 238898 533125 239134
rect 532805 238866 533125 238898
rect 554874 239454 555194 239486
rect 554874 239218 554916 239454
rect 555152 239218 555194 239454
rect 554874 239134 555194 239218
rect 554874 238898 554916 239134
rect 555152 238898 555194 239134
rect 554874 238866 555194 238898
rect 560805 239454 561125 239486
rect 560805 239218 560847 239454
rect 561083 239218 561125 239454
rect 560805 239134 561125 239218
rect 560805 238898 560847 239134
rect 561083 238898 561125 239134
rect 560805 238866 561125 238898
rect -2006 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 -1386 215829
rect -2006 215509 -1386 215593
rect -2006 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 -1386 215509
rect -2006 188829 -1386 215273
rect 19910 215829 20230 215861
rect 19910 215593 19952 215829
rect 20188 215593 20230 215829
rect 19910 215509 20230 215593
rect 19910 215273 19952 215509
rect 20188 215273 20230 215509
rect 19910 215241 20230 215273
rect 25840 215829 26160 215861
rect 25840 215593 25882 215829
rect 26118 215593 26160 215829
rect 25840 215509 26160 215593
rect 25840 215273 25882 215509
rect 26118 215273 26160 215509
rect 25840 215241 26160 215273
rect 31771 215829 32091 215861
rect 31771 215593 31813 215829
rect 32049 215593 32091 215829
rect 31771 215509 32091 215593
rect 31771 215273 31813 215509
rect 32049 215273 32091 215509
rect 31771 215241 32091 215273
rect 47910 215829 48230 215861
rect 47910 215593 47952 215829
rect 48188 215593 48230 215829
rect 47910 215509 48230 215593
rect 47910 215273 47952 215509
rect 48188 215273 48230 215509
rect 47910 215241 48230 215273
rect 53840 215829 54160 215861
rect 53840 215593 53882 215829
rect 54118 215593 54160 215829
rect 53840 215509 54160 215593
rect 53840 215273 53882 215509
rect 54118 215273 54160 215509
rect 53840 215241 54160 215273
rect 59771 215829 60091 215861
rect 59771 215593 59813 215829
rect 60049 215593 60091 215829
rect 59771 215509 60091 215593
rect 59771 215273 59813 215509
rect 60049 215273 60091 215509
rect 59771 215241 60091 215273
rect 75910 215829 76230 215861
rect 75910 215593 75952 215829
rect 76188 215593 76230 215829
rect 75910 215509 76230 215593
rect 75910 215273 75952 215509
rect 76188 215273 76230 215509
rect 75910 215241 76230 215273
rect 81840 215829 82160 215861
rect 81840 215593 81882 215829
rect 82118 215593 82160 215829
rect 81840 215509 82160 215593
rect 81840 215273 81882 215509
rect 82118 215273 82160 215509
rect 81840 215241 82160 215273
rect 87771 215829 88091 215861
rect 87771 215593 87813 215829
rect 88049 215593 88091 215829
rect 87771 215509 88091 215593
rect 87771 215273 87813 215509
rect 88049 215273 88091 215509
rect 87771 215241 88091 215273
rect 103910 215829 104230 215861
rect 103910 215593 103952 215829
rect 104188 215593 104230 215829
rect 103910 215509 104230 215593
rect 103910 215273 103952 215509
rect 104188 215273 104230 215509
rect 103910 215241 104230 215273
rect 109840 215829 110160 215861
rect 109840 215593 109882 215829
rect 110118 215593 110160 215829
rect 109840 215509 110160 215593
rect 109840 215273 109882 215509
rect 110118 215273 110160 215509
rect 109840 215241 110160 215273
rect 115771 215829 116091 215861
rect 115771 215593 115813 215829
rect 116049 215593 116091 215829
rect 115771 215509 116091 215593
rect 115771 215273 115813 215509
rect 116049 215273 116091 215509
rect 115771 215241 116091 215273
rect 131910 215829 132230 215861
rect 131910 215593 131952 215829
rect 132188 215593 132230 215829
rect 131910 215509 132230 215593
rect 131910 215273 131952 215509
rect 132188 215273 132230 215509
rect 131910 215241 132230 215273
rect 137840 215829 138160 215861
rect 137840 215593 137882 215829
rect 138118 215593 138160 215829
rect 137840 215509 138160 215593
rect 137840 215273 137882 215509
rect 138118 215273 138160 215509
rect 137840 215241 138160 215273
rect 143771 215829 144091 215861
rect 143771 215593 143813 215829
rect 144049 215593 144091 215829
rect 143771 215509 144091 215593
rect 143771 215273 143813 215509
rect 144049 215273 144091 215509
rect 143771 215241 144091 215273
rect 159910 215829 160230 215861
rect 159910 215593 159952 215829
rect 160188 215593 160230 215829
rect 159910 215509 160230 215593
rect 159910 215273 159952 215509
rect 160188 215273 160230 215509
rect 159910 215241 160230 215273
rect 165840 215829 166160 215861
rect 165840 215593 165882 215829
rect 166118 215593 166160 215829
rect 165840 215509 166160 215593
rect 165840 215273 165882 215509
rect 166118 215273 166160 215509
rect 165840 215241 166160 215273
rect 171771 215829 172091 215861
rect 171771 215593 171813 215829
rect 172049 215593 172091 215829
rect 171771 215509 172091 215593
rect 171771 215273 171813 215509
rect 172049 215273 172091 215509
rect 171771 215241 172091 215273
rect 187910 215829 188230 215861
rect 187910 215593 187952 215829
rect 188188 215593 188230 215829
rect 187910 215509 188230 215593
rect 187910 215273 187952 215509
rect 188188 215273 188230 215509
rect 187910 215241 188230 215273
rect 193840 215829 194160 215861
rect 193840 215593 193882 215829
rect 194118 215593 194160 215829
rect 193840 215509 194160 215593
rect 193840 215273 193882 215509
rect 194118 215273 194160 215509
rect 193840 215241 194160 215273
rect 199771 215829 200091 215861
rect 199771 215593 199813 215829
rect 200049 215593 200091 215829
rect 199771 215509 200091 215593
rect 199771 215273 199813 215509
rect 200049 215273 200091 215509
rect 199771 215241 200091 215273
rect 215910 215829 216230 215861
rect 215910 215593 215952 215829
rect 216188 215593 216230 215829
rect 215910 215509 216230 215593
rect 215910 215273 215952 215509
rect 216188 215273 216230 215509
rect 215910 215241 216230 215273
rect 221840 215829 222160 215861
rect 221840 215593 221882 215829
rect 222118 215593 222160 215829
rect 221840 215509 222160 215593
rect 221840 215273 221882 215509
rect 222118 215273 222160 215509
rect 221840 215241 222160 215273
rect 227771 215829 228091 215861
rect 227771 215593 227813 215829
rect 228049 215593 228091 215829
rect 227771 215509 228091 215593
rect 227771 215273 227813 215509
rect 228049 215273 228091 215509
rect 227771 215241 228091 215273
rect 243910 215829 244230 215861
rect 243910 215593 243952 215829
rect 244188 215593 244230 215829
rect 243910 215509 244230 215593
rect 243910 215273 243952 215509
rect 244188 215273 244230 215509
rect 243910 215241 244230 215273
rect 249840 215829 250160 215861
rect 249840 215593 249882 215829
rect 250118 215593 250160 215829
rect 249840 215509 250160 215593
rect 249840 215273 249882 215509
rect 250118 215273 250160 215509
rect 249840 215241 250160 215273
rect 255771 215829 256091 215861
rect 255771 215593 255813 215829
rect 256049 215593 256091 215829
rect 255771 215509 256091 215593
rect 255771 215273 255813 215509
rect 256049 215273 256091 215509
rect 255771 215241 256091 215273
rect 271910 215829 272230 215861
rect 271910 215593 271952 215829
rect 272188 215593 272230 215829
rect 271910 215509 272230 215593
rect 271910 215273 271952 215509
rect 272188 215273 272230 215509
rect 271910 215241 272230 215273
rect 277840 215829 278160 215861
rect 277840 215593 277882 215829
rect 278118 215593 278160 215829
rect 277840 215509 278160 215593
rect 277840 215273 277882 215509
rect 278118 215273 278160 215509
rect 277840 215241 278160 215273
rect 283771 215829 284091 215861
rect 283771 215593 283813 215829
rect 284049 215593 284091 215829
rect 283771 215509 284091 215593
rect 283771 215273 283813 215509
rect 284049 215273 284091 215509
rect 283771 215241 284091 215273
rect 299910 215829 300230 215861
rect 299910 215593 299952 215829
rect 300188 215593 300230 215829
rect 299910 215509 300230 215593
rect 299910 215273 299952 215509
rect 300188 215273 300230 215509
rect 299910 215241 300230 215273
rect 305840 215829 306160 215861
rect 305840 215593 305882 215829
rect 306118 215593 306160 215829
rect 305840 215509 306160 215593
rect 305840 215273 305882 215509
rect 306118 215273 306160 215509
rect 305840 215241 306160 215273
rect 311771 215829 312091 215861
rect 311771 215593 311813 215829
rect 312049 215593 312091 215829
rect 311771 215509 312091 215593
rect 311771 215273 311813 215509
rect 312049 215273 312091 215509
rect 311771 215241 312091 215273
rect 327910 215829 328230 215861
rect 327910 215593 327952 215829
rect 328188 215593 328230 215829
rect 327910 215509 328230 215593
rect 327910 215273 327952 215509
rect 328188 215273 328230 215509
rect 327910 215241 328230 215273
rect 333840 215829 334160 215861
rect 333840 215593 333882 215829
rect 334118 215593 334160 215829
rect 333840 215509 334160 215593
rect 333840 215273 333882 215509
rect 334118 215273 334160 215509
rect 333840 215241 334160 215273
rect 339771 215829 340091 215861
rect 339771 215593 339813 215829
rect 340049 215593 340091 215829
rect 339771 215509 340091 215593
rect 339771 215273 339813 215509
rect 340049 215273 340091 215509
rect 339771 215241 340091 215273
rect 355910 215829 356230 215861
rect 355910 215593 355952 215829
rect 356188 215593 356230 215829
rect 355910 215509 356230 215593
rect 355910 215273 355952 215509
rect 356188 215273 356230 215509
rect 355910 215241 356230 215273
rect 361840 215829 362160 215861
rect 361840 215593 361882 215829
rect 362118 215593 362160 215829
rect 361840 215509 362160 215593
rect 361840 215273 361882 215509
rect 362118 215273 362160 215509
rect 361840 215241 362160 215273
rect 367771 215829 368091 215861
rect 367771 215593 367813 215829
rect 368049 215593 368091 215829
rect 367771 215509 368091 215593
rect 367771 215273 367813 215509
rect 368049 215273 368091 215509
rect 367771 215241 368091 215273
rect 383910 215829 384230 215861
rect 383910 215593 383952 215829
rect 384188 215593 384230 215829
rect 383910 215509 384230 215593
rect 383910 215273 383952 215509
rect 384188 215273 384230 215509
rect 383910 215241 384230 215273
rect 389840 215829 390160 215861
rect 389840 215593 389882 215829
rect 390118 215593 390160 215829
rect 389840 215509 390160 215593
rect 389840 215273 389882 215509
rect 390118 215273 390160 215509
rect 389840 215241 390160 215273
rect 395771 215829 396091 215861
rect 395771 215593 395813 215829
rect 396049 215593 396091 215829
rect 395771 215509 396091 215593
rect 395771 215273 395813 215509
rect 396049 215273 396091 215509
rect 395771 215241 396091 215273
rect 411910 215829 412230 215861
rect 411910 215593 411952 215829
rect 412188 215593 412230 215829
rect 411910 215509 412230 215593
rect 411910 215273 411952 215509
rect 412188 215273 412230 215509
rect 411910 215241 412230 215273
rect 417840 215829 418160 215861
rect 417840 215593 417882 215829
rect 418118 215593 418160 215829
rect 417840 215509 418160 215593
rect 417840 215273 417882 215509
rect 418118 215273 418160 215509
rect 417840 215241 418160 215273
rect 423771 215829 424091 215861
rect 423771 215593 423813 215829
rect 424049 215593 424091 215829
rect 423771 215509 424091 215593
rect 423771 215273 423813 215509
rect 424049 215273 424091 215509
rect 423771 215241 424091 215273
rect 439910 215829 440230 215861
rect 439910 215593 439952 215829
rect 440188 215593 440230 215829
rect 439910 215509 440230 215593
rect 439910 215273 439952 215509
rect 440188 215273 440230 215509
rect 439910 215241 440230 215273
rect 445840 215829 446160 215861
rect 445840 215593 445882 215829
rect 446118 215593 446160 215829
rect 445840 215509 446160 215593
rect 445840 215273 445882 215509
rect 446118 215273 446160 215509
rect 445840 215241 446160 215273
rect 451771 215829 452091 215861
rect 451771 215593 451813 215829
rect 452049 215593 452091 215829
rect 451771 215509 452091 215593
rect 451771 215273 451813 215509
rect 452049 215273 452091 215509
rect 451771 215241 452091 215273
rect 467910 215829 468230 215861
rect 467910 215593 467952 215829
rect 468188 215593 468230 215829
rect 467910 215509 468230 215593
rect 467910 215273 467952 215509
rect 468188 215273 468230 215509
rect 467910 215241 468230 215273
rect 473840 215829 474160 215861
rect 473840 215593 473882 215829
rect 474118 215593 474160 215829
rect 473840 215509 474160 215593
rect 473840 215273 473882 215509
rect 474118 215273 474160 215509
rect 473840 215241 474160 215273
rect 479771 215829 480091 215861
rect 479771 215593 479813 215829
rect 480049 215593 480091 215829
rect 479771 215509 480091 215593
rect 479771 215273 479813 215509
rect 480049 215273 480091 215509
rect 479771 215241 480091 215273
rect 495910 215829 496230 215861
rect 495910 215593 495952 215829
rect 496188 215593 496230 215829
rect 495910 215509 496230 215593
rect 495910 215273 495952 215509
rect 496188 215273 496230 215509
rect 495910 215241 496230 215273
rect 501840 215829 502160 215861
rect 501840 215593 501882 215829
rect 502118 215593 502160 215829
rect 501840 215509 502160 215593
rect 501840 215273 501882 215509
rect 502118 215273 502160 215509
rect 501840 215241 502160 215273
rect 507771 215829 508091 215861
rect 507771 215593 507813 215829
rect 508049 215593 508091 215829
rect 507771 215509 508091 215593
rect 507771 215273 507813 215509
rect 508049 215273 508091 215509
rect 507771 215241 508091 215273
rect 523910 215829 524230 215861
rect 523910 215593 523952 215829
rect 524188 215593 524230 215829
rect 523910 215509 524230 215593
rect 523910 215273 523952 215509
rect 524188 215273 524230 215509
rect 523910 215241 524230 215273
rect 529840 215829 530160 215861
rect 529840 215593 529882 215829
rect 530118 215593 530160 215829
rect 529840 215509 530160 215593
rect 529840 215273 529882 215509
rect 530118 215273 530160 215509
rect 529840 215241 530160 215273
rect 535771 215829 536091 215861
rect 535771 215593 535813 215829
rect 536049 215593 536091 215829
rect 535771 215509 536091 215593
rect 535771 215273 535813 215509
rect 536049 215273 536091 215509
rect 535771 215241 536091 215273
rect 551910 215829 552230 215861
rect 551910 215593 551952 215829
rect 552188 215593 552230 215829
rect 551910 215509 552230 215593
rect 551910 215273 551952 215509
rect 552188 215273 552230 215509
rect 551910 215241 552230 215273
rect 557840 215829 558160 215861
rect 557840 215593 557882 215829
rect 558118 215593 558160 215829
rect 557840 215509 558160 215593
rect 557840 215273 557882 215509
rect 558118 215273 558160 215509
rect 557840 215241 558160 215273
rect 563771 215829 564091 215861
rect 563771 215593 563813 215829
rect 564049 215593 564091 215829
rect 563771 215509 564091 215593
rect 563771 215273 563813 215509
rect 564049 215273 564091 215509
rect 563771 215241 564091 215273
rect 573494 215829 574114 242273
rect 573494 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 574114 215829
rect 573494 215509 574114 215593
rect 573494 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 574114 215509
rect 22874 212454 23194 212486
rect 22874 212218 22916 212454
rect 23152 212218 23194 212454
rect 22874 212134 23194 212218
rect 22874 211898 22916 212134
rect 23152 211898 23194 212134
rect 22874 211866 23194 211898
rect 28805 212454 29125 212486
rect 28805 212218 28847 212454
rect 29083 212218 29125 212454
rect 28805 212134 29125 212218
rect 28805 211898 28847 212134
rect 29083 211898 29125 212134
rect 28805 211866 29125 211898
rect 50874 212454 51194 212486
rect 50874 212218 50916 212454
rect 51152 212218 51194 212454
rect 50874 212134 51194 212218
rect 50874 211898 50916 212134
rect 51152 211898 51194 212134
rect 50874 211866 51194 211898
rect 56805 212454 57125 212486
rect 56805 212218 56847 212454
rect 57083 212218 57125 212454
rect 56805 212134 57125 212218
rect 56805 211898 56847 212134
rect 57083 211898 57125 212134
rect 56805 211866 57125 211898
rect 78874 212454 79194 212486
rect 78874 212218 78916 212454
rect 79152 212218 79194 212454
rect 78874 212134 79194 212218
rect 78874 211898 78916 212134
rect 79152 211898 79194 212134
rect 78874 211866 79194 211898
rect 84805 212454 85125 212486
rect 84805 212218 84847 212454
rect 85083 212218 85125 212454
rect 84805 212134 85125 212218
rect 84805 211898 84847 212134
rect 85083 211898 85125 212134
rect 84805 211866 85125 211898
rect 106874 212454 107194 212486
rect 106874 212218 106916 212454
rect 107152 212218 107194 212454
rect 106874 212134 107194 212218
rect 106874 211898 106916 212134
rect 107152 211898 107194 212134
rect 106874 211866 107194 211898
rect 112805 212454 113125 212486
rect 112805 212218 112847 212454
rect 113083 212218 113125 212454
rect 112805 212134 113125 212218
rect 112805 211898 112847 212134
rect 113083 211898 113125 212134
rect 112805 211866 113125 211898
rect 134874 212454 135194 212486
rect 134874 212218 134916 212454
rect 135152 212218 135194 212454
rect 134874 212134 135194 212218
rect 134874 211898 134916 212134
rect 135152 211898 135194 212134
rect 134874 211866 135194 211898
rect 140805 212454 141125 212486
rect 140805 212218 140847 212454
rect 141083 212218 141125 212454
rect 140805 212134 141125 212218
rect 140805 211898 140847 212134
rect 141083 211898 141125 212134
rect 140805 211866 141125 211898
rect 162874 212454 163194 212486
rect 162874 212218 162916 212454
rect 163152 212218 163194 212454
rect 162874 212134 163194 212218
rect 162874 211898 162916 212134
rect 163152 211898 163194 212134
rect 162874 211866 163194 211898
rect 168805 212454 169125 212486
rect 168805 212218 168847 212454
rect 169083 212218 169125 212454
rect 168805 212134 169125 212218
rect 168805 211898 168847 212134
rect 169083 211898 169125 212134
rect 168805 211866 169125 211898
rect 190874 212454 191194 212486
rect 190874 212218 190916 212454
rect 191152 212218 191194 212454
rect 190874 212134 191194 212218
rect 190874 211898 190916 212134
rect 191152 211898 191194 212134
rect 190874 211866 191194 211898
rect 196805 212454 197125 212486
rect 196805 212218 196847 212454
rect 197083 212218 197125 212454
rect 196805 212134 197125 212218
rect 196805 211898 196847 212134
rect 197083 211898 197125 212134
rect 196805 211866 197125 211898
rect 218874 212454 219194 212486
rect 218874 212218 218916 212454
rect 219152 212218 219194 212454
rect 218874 212134 219194 212218
rect 218874 211898 218916 212134
rect 219152 211898 219194 212134
rect 218874 211866 219194 211898
rect 224805 212454 225125 212486
rect 224805 212218 224847 212454
rect 225083 212218 225125 212454
rect 224805 212134 225125 212218
rect 224805 211898 224847 212134
rect 225083 211898 225125 212134
rect 224805 211866 225125 211898
rect 246874 212454 247194 212486
rect 246874 212218 246916 212454
rect 247152 212218 247194 212454
rect 246874 212134 247194 212218
rect 246874 211898 246916 212134
rect 247152 211898 247194 212134
rect 246874 211866 247194 211898
rect 252805 212454 253125 212486
rect 252805 212218 252847 212454
rect 253083 212218 253125 212454
rect 252805 212134 253125 212218
rect 252805 211898 252847 212134
rect 253083 211898 253125 212134
rect 252805 211866 253125 211898
rect 274874 212454 275194 212486
rect 274874 212218 274916 212454
rect 275152 212218 275194 212454
rect 274874 212134 275194 212218
rect 274874 211898 274916 212134
rect 275152 211898 275194 212134
rect 274874 211866 275194 211898
rect 280805 212454 281125 212486
rect 280805 212218 280847 212454
rect 281083 212218 281125 212454
rect 280805 212134 281125 212218
rect 280805 211898 280847 212134
rect 281083 211898 281125 212134
rect 280805 211866 281125 211898
rect 302874 212454 303194 212486
rect 302874 212218 302916 212454
rect 303152 212218 303194 212454
rect 302874 212134 303194 212218
rect 302874 211898 302916 212134
rect 303152 211898 303194 212134
rect 302874 211866 303194 211898
rect 308805 212454 309125 212486
rect 308805 212218 308847 212454
rect 309083 212218 309125 212454
rect 308805 212134 309125 212218
rect 308805 211898 308847 212134
rect 309083 211898 309125 212134
rect 308805 211866 309125 211898
rect 330874 212454 331194 212486
rect 330874 212218 330916 212454
rect 331152 212218 331194 212454
rect 330874 212134 331194 212218
rect 330874 211898 330916 212134
rect 331152 211898 331194 212134
rect 330874 211866 331194 211898
rect 336805 212454 337125 212486
rect 336805 212218 336847 212454
rect 337083 212218 337125 212454
rect 336805 212134 337125 212218
rect 336805 211898 336847 212134
rect 337083 211898 337125 212134
rect 336805 211866 337125 211898
rect 358874 212454 359194 212486
rect 358874 212218 358916 212454
rect 359152 212218 359194 212454
rect 358874 212134 359194 212218
rect 358874 211898 358916 212134
rect 359152 211898 359194 212134
rect 358874 211866 359194 211898
rect 364805 212454 365125 212486
rect 364805 212218 364847 212454
rect 365083 212218 365125 212454
rect 364805 212134 365125 212218
rect 364805 211898 364847 212134
rect 365083 211898 365125 212134
rect 364805 211866 365125 211898
rect 386874 212454 387194 212486
rect 386874 212218 386916 212454
rect 387152 212218 387194 212454
rect 386874 212134 387194 212218
rect 386874 211898 386916 212134
rect 387152 211898 387194 212134
rect 386874 211866 387194 211898
rect 392805 212454 393125 212486
rect 392805 212218 392847 212454
rect 393083 212218 393125 212454
rect 392805 212134 393125 212218
rect 392805 211898 392847 212134
rect 393083 211898 393125 212134
rect 392805 211866 393125 211898
rect 414874 212454 415194 212486
rect 414874 212218 414916 212454
rect 415152 212218 415194 212454
rect 414874 212134 415194 212218
rect 414874 211898 414916 212134
rect 415152 211898 415194 212134
rect 414874 211866 415194 211898
rect 420805 212454 421125 212486
rect 420805 212218 420847 212454
rect 421083 212218 421125 212454
rect 420805 212134 421125 212218
rect 420805 211898 420847 212134
rect 421083 211898 421125 212134
rect 420805 211866 421125 211898
rect 442874 212454 443194 212486
rect 442874 212218 442916 212454
rect 443152 212218 443194 212454
rect 442874 212134 443194 212218
rect 442874 211898 442916 212134
rect 443152 211898 443194 212134
rect 442874 211866 443194 211898
rect 448805 212454 449125 212486
rect 448805 212218 448847 212454
rect 449083 212218 449125 212454
rect 448805 212134 449125 212218
rect 448805 211898 448847 212134
rect 449083 211898 449125 212134
rect 448805 211866 449125 211898
rect 470874 212454 471194 212486
rect 470874 212218 470916 212454
rect 471152 212218 471194 212454
rect 470874 212134 471194 212218
rect 470874 211898 470916 212134
rect 471152 211898 471194 212134
rect 470874 211866 471194 211898
rect 476805 212454 477125 212486
rect 476805 212218 476847 212454
rect 477083 212218 477125 212454
rect 476805 212134 477125 212218
rect 476805 211898 476847 212134
rect 477083 211898 477125 212134
rect 476805 211866 477125 211898
rect 498874 212454 499194 212486
rect 498874 212218 498916 212454
rect 499152 212218 499194 212454
rect 498874 212134 499194 212218
rect 498874 211898 498916 212134
rect 499152 211898 499194 212134
rect 498874 211866 499194 211898
rect 504805 212454 505125 212486
rect 504805 212218 504847 212454
rect 505083 212218 505125 212454
rect 504805 212134 505125 212218
rect 504805 211898 504847 212134
rect 505083 211898 505125 212134
rect 504805 211866 505125 211898
rect 526874 212454 527194 212486
rect 526874 212218 526916 212454
rect 527152 212218 527194 212454
rect 526874 212134 527194 212218
rect 526874 211898 526916 212134
rect 527152 211898 527194 212134
rect 526874 211866 527194 211898
rect 532805 212454 533125 212486
rect 532805 212218 532847 212454
rect 533083 212218 533125 212454
rect 532805 212134 533125 212218
rect 532805 211898 532847 212134
rect 533083 211898 533125 212134
rect 532805 211866 533125 211898
rect 554874 212454 555194 212486
rect 554874 212218 554916 212454
rect 555152 212218 555194 212454
rect 554874 212134 555194 212218
rect 554874 211898 554916 212134
rect 555152 211898 555194 212134
rect 554874 211866 555194 211898
rect 560805 212454 561125 212486
rect 560805 212218 560847 212454
rect 561083 212218 561125 212454
rect 560805 212134 561125 212218
rect 560805 211898 560847 212134
rect 561083 211898 561125 212134
rect 560805 211866 561125 211898
rect -2006 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 -1386 188829
rect -2006 188509 -1386 188593
rect -2006 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 -1386 188509
rect -2006 161829 -1386 188273
rect 19910 188829 20230 188861
rect 19910 188593 19952 188829
rect 20188 188593 20230 188829
rect 19910 188509 20230 188593
rect 19910 188273 19952 188509
rect 20188 188273 20230 188509
rect 19910 188241 20230 188273
rect 25840 188829 26160 188861
rect 25840 188593 25882 188829
rect 26118 188593 26160 188829
rect 25840 188509 26160 188593
rect 25840 188273 25882 188509
rect 26118 188273 26160 188509
rect 25840 188241 26160 188273
rect 31771 188829 32091 188861
rect 31771 188593 31813 188829
rect 32049 188593 32091 188829
rect 31771 188509 32091 188593
rect 31771 188273 31813 188509
rect 32049 188273 32091 188509
rect 31771 188241 32091 188273
rect 47910 188829 48230 188861
rect 47910 188593 47952 188829
rect 48188 188593 48230 188829
rect 47910 188509 48230 188593
rect 47910 188273 47952 188509
rect 48188 188273 48230 188509
rect 47910 188241 48230 188273
rect 53840 188829 54160 188861
rect 53840 188593 53882 188829
rect 54118 188593 54160 188829
rect 53840 188509 54160 188593
rect 53840 188273 53882 188509
rect 54118 188273 54160 188509
rect 53840 188241 54160 188273
rect 59771 188829 60091 188861
rect 59771 188593 59813 188829
rect 60049 188593 60091 188829
rect 59771 188509 60091 188593
rect 59771 188273 59813 188509
rect 60049 188273 60091 188509
rect 59771 188241 60091 188273
rect 75910 188829 76230 188861
rect 75910 188593 75952 188829
rect 76188 188593 76230 188829
rect 75910 188509 76230 188593
rect 75910 188273 75952 188509
rect 76188 188273 76230 188509
rect 75910 188241 76230 188273
rect 81840 188829 82160 188861
rect 81840 188593 81882 188829
rect 82118 188593 82160 188829
rect 81840 188509 82160 188593
rect 81840 188273 81882 188509
rect 82118 188273 82160 188509
rect 81840 188241 82160 188273
rect 87771 188829 88091 188861
rect 87771 188593 87813 188829
rect 88049 188593 88091 188829
rect 87771 188509 88091 188593
rect 87771 188273 87813 188509
rect 88049 188273 88091 188509
rect 87771 188241 88091 188273
rect 103910 188829 104230 188861
rect 103910 188593 103952 188829
rect 104188 188593 104230 188829
rect 103910 188509 104230 188593
rect 103910 188273 103952 188509
rect 104188 188273 104230 188509
rect 103910 188241 104230 188273
rect 109840 188829 110160 188861
rect 109840 188593 109882 188829
rect 110118 188593 110160 188829
rect 109840 188509 110160 188593
rect 109840 188273 109882 188509
rect 110118 188273 110160 188509
rect 109840 188241 110160 188273
rect 115771 188829 116091 188861
rect 115771 188593 115813 188829
rect 116049 188593 116091 188829
rect 115771 188509 116091 188593
rect 115771 188273 115813 188509
rect 116049 188273 116091 188509
rect 115771 188241 116091 188273
rect 131910 188829 132230 188861
rect 131910 188593 131952 188829
rect 132188 188593 132230 188829
rect 131910 188509 132230 188593
rect 131910 188273 131952 188509
rect 132188 188273 132230 188509
rect 131910 188241 132230 188273
rect 137840 188829 138160 188861
rect 137840 188593 137882 188829
rect 138118 188593 138160 188829
rect 137840 188509 138160 188593
rect 137840 188273 137882 188509
rect 138118 188273 138160 188509
rect 137840 188241 138160 188273
rect 143771 188829 144091 188861
rect 143771 188593 143813 188829
rect 144049 188593 144091 188829
rect 143771 188509 144091 188593
rect 143771 188273 143813 188509
rect 144049 188273 144091 188509
rect 143771 188241 144091 188273
rect 159910 188829 160230 188861
rect 159910 188593 159952 188829
rect 160188 188593 160230 188829
rect 159910 188509 160230 188593
rect 159910 188273 159952 188509
rect 160188 188273 160230 188509
rect 159910 188241 160230 188273
rect 165840 188829 166160 188861
rect 165840 188593 165882 188829
rect 166118 188593 166160 188829
rect 165840 188509 166160 188593
rect 165840 188273 165882 188509
rect 166118 188273 166160 188509
rect 165840 188241 166160 188273
rect 171771 188829 172091 188861
rect 171771 188593 171813 188829
rect 172049 188593 172091 188829
rect 171771 188509 172091 188593
rect 171771 188273 171813 188509
rect 172049 188273 172091 188509
rect 171771 188241 172091 188273
rect 187910 188829 188230 188861
rect 187910 188593 187952 188829
rect 188188 188593 188230 188829
rect 187910 188509 188230 188593
rect 187910 188273 187952 188509
rect 188188 188273 188230 188509
rect 187910 188241 188230 188273
rect 193840 188829 194160 188861
rect 193840 188593 193882 188829
rect 194118 188593 194160 188829
rect 193840 188509 194160 188593
rect 193840 188273 193882 188509
rect 194118 188273 194160 188509
rect 193840 188241 194160 188273
rect 199771 188829 200091 188861
rect 199771 188593 199813 188829
rect 200049 188593 200091 188829
rect 199771 188509 200091 188593
rect 199771 188273 199813 188509
rect 200049 188273 200091 188509
rect 199771 188241 200091 188273
rect 215910 188829 216230 188861
rect 215910 188593 215952 188829
rect 216188 188593 216230 188829
rect 215910 188509 216230 188593
rect 215910 188273 215952 188509
rect 216188 188273 216230 188509
rect 215910 188241 216230 188273
rect 221840 188829 222160 188861
rect 221840 188593 221882 188829
rect 222118 188593 222160 188829
rect 221840 188509 222160 188593
rect 221840 188273 221882 188509
rect 222118 188273 222160 188509
rect 221840 188241 222160 188273
rect 227771 188829 228091 188861
rect 227771 188593 227813 188829
rect 228049 188593 228091 188829
rect 227771 188509 228091 188593
rect 227771 188273 227813 188509
rect 228049 188273 228091 188509
rect 227771 188241 228091 188273
rect 243910 188829 244230 188861
rect 243910 188593 243952 188829
rect 244188 188593 244230 188829
rect 243910 188509 244230 188593
rect 243910 188273 243952 188509
rect 244188 188273 244230 188509
rect 243910 188241 244230 188273
rect 249840 188829 250160 188861
rect 249840 188593 249882 188829
rect 250118 188593 250160 188829
rect 249840 188509 250160 188593
rect 249840 188273 249882 188509
rect 250118 188273 250160 188509
rect 249840 188241 250160 188273
rect 255771 188829 256091 188861
rect 255771 188593 255813 188829
rect 256049 188593 256091 188829
rect 255771 188509 256091 188593
rect 255771 188273 255813 188509
rect 256049 188273 256091 188509
rect 255771 188241 256091 188273
rect 271910 188829 272230 188861
rect 271910 188593 271952 188829
rect 272188 188593 272230 188829
rect 271910 188509 272230 188593
rect 271910 188273 271952 188509
rect 272188 188273 272230 188509
rect 271910 188241 272230 188273
rect 277840 188829 278160 188861
rect 277840 188593 277882 188829
rect 278118 188593 278160 188829
rect 277840 188509 278160 188593
rect 277840 188273 277882 188509
rect 278118 188273 278160 188509
rect 277840 188241 278160 188273
rect 283771 188829 284091 188861
rect 283771 188593 283813 188829
rect 284049 188593 284091 188829
rect 283771 188509 284091 188593
rect 283771 188273 283813 188509
rect 284049 188273 284091 188509
rect 283771 188241 284091 188273
rect 299910 188829 300230 188861
rect 299910 188593 299952 188829
rect 300188 188593 300230 188829
rect 299910 188509 300230 188593
rect 299910 188273 299952 188509
rect 300188 188273 300230 188509
rect 299910 188241 300230 188273
rect 305840 188829 306160 188861
rect 305840 188593 305882 188829
rect 306118 188593 306160 188829
rect 305840 188509 306160 188593
rect 305840 188273 305882 188509
rect 306118 188273 306160 188509
rect 305840 188241 306160 188273
rect 311771 188829 312091 188861
rect 311771 188593 311813 188829
rect 312049 188593 312091 188829
rect 311771 188509 312091 188593
rect 311771 188273 311813 188509
rect 312049 188273 312091 188509
rect 311771 188241 312091 188273
rect 327910 188829 328230 188861
rect 327910 188593 327952 188829
rect 328188 188593 328230 188829
rect 327910 188509 328230 188593
rect 327910 188273 327952 188509
rect 328188 188273 328230 188509
rect 327910 188241 328230 188273
rect 333840 188829 334160 188861
rect 333840 188593 333882 188829
rect 334118 188593 334160 188829
rect 333840 188509 334160 188593
rect 333840 188273 333882 188509
rect 334118 188273 334160 188509
rect 333840 188241 334160 188273
rect 339771 188829 340091 188861
rect 339771 188593 339813 188829
rect 340049 188593 340091 188829
rect 339771 188509 340091 188593
rect 339771 188273 339813 188509
rect 340049 188273 340091 188509
rect 339771 188241 340091 188273
rect 355910 188829 356230 188861
rect 355910 188593 355952 188829
rect 356188 188593 356230 188829
rect 355910 188509 356230 188593
rect 355910 188273 355952 188509
rect 356188 188273 356230 188509
rect 355910 188241 356230 188273
rect 361840 188829 362160 188861
rect 361840 188593 361882 188829
rect 362118 188593 362160 188829
rect 361840 188509 362160 188593
rect 361840 188273 361882 188509
rect 362118 188273 362160 188509
rect 361840 188241 362160 188273
rect 367771 188829 368091 188861
rect 367771 188593 367813 188829
rect 368049 188593 368091 188829
rect 367771 188509 368091 188593
rect 367771 188273 367813 188509
rect 368049 188273 368091 188509
rect 367771 188241 368091 188273
rect 383910 188829 384230 188861
rect 383910 188593 383952 188829
rect 384188 188593 384230 188829
rect 383910 188509 384230 188593
rect 383910 188273 383952 188509
rect 384188 188273 384230 188509
rect 383910 188241 384230 188273
rect 389840 188829 390160 188861
rect 389840 188593 389882 188829
rect 390118 188593 390160 188829
rect 389840 188509 390160 188593
rect 389840 188273 389882 188509
rect 390118 188273 390160 188509
rect 389840 188241 390160 188273
rect 395771 188829 396091 188861
rect 395771 188593 395813 188829
rect 396049 188593 396091 188829
rect 395771 188509 396091 188593
rect 395771 188273 395813 188509
rect 396049 188273 396091 188509
rect 395771 188241 396091 188273
rect 411910 188829 412230 188861
rect 411910 188593 411952 188829
rect 412188 188593 412230 188829
rect 411910 188509 412230 188593
rect 411910 188273 411952 188509
rect 412188 188273 412230 188509
rect 411910 188241 412230 188273
rect 417840 188829 418160 188861
rect 417840 188593 417882 188829
rect 418118 188593 418160 188829
rect 417840 188509 418160 188593
rect 417840 188273 417882 188509
rect 418118 188273 418160 188509
rect 417840 188241 418160 188273
rect 423771 188829 424091 188861
rect 423771 188593 423813 188829
rect 424049 188593 424091 188829
rect 423771 188509 424091 188593
rect 423771 188273 423813 188509
rect 424049 188273 424091 188509
rect 423771 188241 424091 188273
rect 439910 188829 440230 188861
rect 439910 188593 439952 188829
rect 440188 188593 440230 188829
rect 439910 188509 440230 188593
rect 439910 188273 439952 188509
rect 440188 188273 440230 188509
rect 439910 188241 440230 188273
rect 445840 188829 446160 188861
rect 445840 188593 445882 188829
rect 446118 188593 446160 188829
rect 445840 188509 446160 188593
rect 445840 188273 445882 188509
rect 446118 188273 446160 188509
rect 445840 188241 446160 188273
rect 451771 188829 452091 188861
rect 451771 188593 451813 188829
rect 452049 188593 452091 188829
rect 451771 188509 452091 188593
rect 451771 188273 451813 188509
rect 452049 188273 452091 188509
rect 451771 188241 452091 188273
rect 467910 188829 468230 188861
rect 467910 188593 467952 188829
rect 468188 188593 468230 188829
rect 467910 188509 468230 188593
rect 467910 188273 467952 188509
rect 468188 188273 468230 188509
rect 467910 188241 468230 188273
rect 473840 188829 474160 188861
rect 473840 188593 473882 188829
rect 474118 188593 474160 188829
rect 473840 188509 474160 188593
rect 473840 188273 473882 188509
rect 474118 188273 474160 188509
rect 473840 188241 474160 188273
rect 479771 188829 480091 188861
rect 479771 188593 479813 188829
rect 480049 188593 480091 188829
rect 479771 188509 480091 188593
rect 479771 188273 479813 188509
rect 480049 188273 480091 188509
rect 479771 188241 480091 188273
rect 495910 188829 496230 188861
rect 495910 188593 495952 188829
rect 496188 188593 496230 188829
rect 495910 188509 496230 188593
rect 495910 188273 495952 188509
rect 496188 188273 496230 188509
rect 495910 188241 496230 188273
rect 501840 188829 502160 188861
rect 501840 188593 501882 188829
rect 502118 188593 502160 188829
rect 501840 188509 502160 188593
rect 501840 188273 501882 188509
rect 502118 188273 502160 188509
rect 501840 188241 502160 188273
rect 507771 188829 508091 188861
rect 507771 188593 507813 188829
rect 508049 188593 508091 188829
rect 507771 188509 508091 188593
rect 507771 188273 507813 188509
rect 508049 188273 508091 188509
rect 507771 188241 508091 188273
rect 523910 188829 524230 188861
rect 523910 188593 523952 188829
rect 524188 188593 524230 188829
rect 523910 188509 524230 188593
rect 523910 188273 523952 188509
rect 524188 188273 524230 188509
rect 523910 188241 524230 188273
rect 529840 188829 530160 188861
rect 529840 188593 529882 188829
rect 530118 188593 530160 188829
rect 529840 188509 530160 188593
rect 529840 188273 529882 188509
rect 530118 188273 530160 188509
rect 529840 188241 530160 188273
rect 535771 188829 536091 188861
rect 535771 188593 535813 188829
rect 536049 188593 536091 188829
rect 535771 188509 536091 188593
rect 535771 188273 535813 188509
rect 536049 188273 536091 188509
rect 535771 188241 536091 188273
rect 551910 188829 552230 188861
rect 551910 188593 551952 188829
rect 552188 188593 552230 188829
rect 551910 188509 552230 188593
rect 551910 188273 551952 188509
rect 552188 188273 552230 188509
rect 551910 188241 552230 188273
rect 557840 188829 558160 188861
rect 557840 188593 557882 188829
rect 558118 188593 558160 188829
rect 557840 188509 558160 188593
rect 557840 188273 557882 188509
rect 558118 188273 558160 188509
rect 557840 188241 558160 188273
rect 563771 188829 564091 188861
rect 563771 188593 563813 188829
rect 564049 188593 564091 188829
rect 563771 188509 564091 188593
rect 563771 188273 563813 188509
rect 564049 188273 564091 188509
rect 563771 188241 564091 188273
rect 573494 188829 574114 215273
rect 573494 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 574114 188829
rect 573494 188509 574114 188593
rect 573494 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 574114 188509
rect 22874 185454 23194 185486
rect 22874 185218 22916 185454
rect 23152 185218 23194 185454
rect 22874 185134 23194 185218
rect 22874 184898 22916 185134
rect 23152 184898 23194 185134
rect 22874 184866 23194 184898
rect 28805 185454 29125 185486
rect 28805 185218 28847 185454
rect 29083 185218 29125 185454
rect 28805 185134 29125 185218
rect 28805 184898 28847 185134
rect 29083 184898 29125 185134
rect 28805 184866 29125 184898
rect 50874 185454 51194 185486
rect 50874 185218 50916 185454
rect 51152 185218 51194 185454
rect 50874 185134 51194 185218
rect 50874 184898 50916 185134
rect 51152 184898 51194 185134
rect 50874 184866 51194 184898
rect 56805 185454 57125 185486
rect 56805 185218 56847 185454
rect 57083 185218 57125 185454
rect 56805 185134 57125 185218
rect 56805 184898 56847 185134
rect 57083 184898 57125 185134
rect 56805 184866 57125 184898
rect 78874 185454 79194 185486
rect 78874 185218 78916 185454
rect 79152 185218 79194 185454
rect 78874 185134 79194 185218
rect 78874 184898 78916 185134
rect 79152 184898 79194 185134
rect 78874 184866 79194 184898
rect 84805 185454 85125 185486
rect 84805 185218 84847 185454
rect 85083 185218 85125 185454
rect 84805 185134 85125 185218
rect 84805 184898 84847 185134
rect 85083 184898 85125 185134
rect 84805 184866 85125 184898
rect 106874 185454 107194 185486
rect 106874 185218 106916 185454
rect 107152 185218 107194 185454
rect 106874 185134 107194 185218
rect 106874 184898 106916 185134
rect 107152 184898 107194 185134
rect 106874 184866 107194 184898
rect 112805 185454 113125 185486
rect 112805 185218 112847 185454
rect 113083 185218 113125 185454
rect 112805 185134 113125 185218
rect 112805 184898 112847 185134
rect 113083 184898 113125 185134
rect 112805 184866 113125 184898
rect 134874 185454 135194 185486
rect 134874 185218 134916 185454
rect 135152 185218 135194 185454
rect 134874 185134 135194 185218
rect 134874 184898 134916 185134
rect 135152 184898 135194 185134
rect 134874 184866 135194 184898
rect 140805 185454 141125 185486
rect 140805 185218 140847 185454
rect 141083 185218 141125 185454
rect 140805 185134 141125 185218
rect 140805 184898 140847 185134
rect 141083 184898 141125 185134
rect 140805 184866 141125 184898
rect 162874 185454 163194 185486
rect 162874 185218 162916 185454
rect 163152 185218 163194 185454
rect 162874 185134 163194 185218
rect 162874 184898 162916 185134
rect 163152 184898 163194 185134
rect 162874 184866 163194 184898
rect 168805 185454 169125 185486
rect 168805 185218 168847 185454
rect 169083 185218 169125 185454
rect 168805 185134 169125 185218
rect 168805 184898 168847 185134
rect 169083 184898 169125 185134
rect 168805 184866 169125 184898
rect 190874 185454 191194 185486
rect 190874 185218 190916 185454
rect 191152 185218 191194 185454
rect 190874 185134 191194 185218
rect 190874 184898 190916 185134
rect 191152 184898 191194 185134
rect 190874 184866 191194 184898
rect 196805 185454 197125 185486
rect 196805 185218 196847 185454
rect 197083 185218 197125 185454
rect 196805 185134 197125 185218
rect 196805 184898 196847 185134
rect 197083 184898 197125 185134
rect 196805 184866 197125 184898
rect 218874 185454 219194 185486
rect 218874 185218 218916 185454
rect 219152 185218 219194 185454
rect 218874 185134 219194 185218
rect 218874 184898 218916 185134
rect 219152 184898 219194 185134
rect 218874 184866 219194 184898
rect 224805 185454 225125 185486
rect 224805 185218 224847 185454
rect 225083 185218 225125 185454
rect 224805 185134 225125 185218
rect 224805 184898 224847 185134
rect 225083 184898 225125 185134
rect 224805 184866 225125 184898
rect 246874 185454 247194 185486
rect 246874 185218 246916 185454
rect 247152 185218 247194 185454
rect 246874 185134 247194 185218
rect 246874 184898 246916 185134
rect 247152 184898 247194 185134
rect 246874 184866 247194 184898
rect 252805 185454 253125 185486
rect 252805 185218 252847 185454
rect 253083 185218 253125 185454
rect 252805 185134 253125 185218
rect 252805 184898 252847 185134
rect 253083 184898 253125 185134
rect 252805 184866 253125 184898
rect 274874 185454 275194 185486
rect 274874 185218 274916 185454
rect 275152 185218 275194 185454
rect 274874 185134 275194 185218
rect 274874 184898 274916 185134
rect 275152 184898 275194 185134
rect 274874 184866 275194 184898
rect 280805 185454 281125 185486
rect 280805 185218 280847 185454
rect 281083 185218 281125 185454
rect 280805 185134 281125 185218
rect 280805 184898 280847 185134
rect 281083 184898 281125 185134
rect 280805 184866 281125 184898
rect 302874 185454 303194 185486
rect 302874 185218 302916 185454
rect 303152 185218 303194 185454
rect 302874 185134 303194 185218
rect 302874 184898 302916 185134
rect 303152 184898 303194 185134
rect 302874 184866 303194 184898
rect 308805 185454 309125 185486
rect 308805 185218 308847 185454
rect 309083 185218 309125 185454
rect 308805 185134 309125 185218
rect 308805 184898 308847 185134
rect 309083 184898 309125 185134
rect 308805 184866 309125 184898
rect 330874 185454 331194 185486
rect 330874 185218 330916 185454
rect 331152 185218 331194 185454
rect 330874 185134 331194 185218
rect 330874 184898 330916 185134
rect 331152 184898 331194 185134
rect 330874 184866 331194 184898
rect 336805 185454 337125 185486
rect 336805 185218 336847 185454
rect 337083 185218 337125 185454
rect 336805 185134 337125 185218
rect 336805 184898 336847 185134
rect 337083 184898 337125 185134
rect 336805 184866 337125 184898
rect 358874 185454 359194 185486
rect 358874 185218 358916 185454
rect 359152 185218 359194 185454
rect 358874 185134 359194 185218
rect 358874 184898 358916 185134
rect 359152 184898 359194 185134
rect 358874 184866 359194 184898
rect 364805 185454 365125 185486
rect 364805 185218 364847 185454
rect 365083 185218 365125 185454
rect 364805 185134 365125 185218
rect 364805 184898 364847 185134
rect 365083 184898 365125 185134
rect 364805 184866 365125 184898
rect 386874 185454 387194 185486
rect 386874 185218 386916 185454
rect 387152 185218 387194 185454
rect 386874 185134 387194 185218
rect 386874 184898 386916 185134
rect 387152 184898 387194 185134
rect 386874 184866 387194 184898
rect 392805 185454 393125 185486
rect 392805 185218 392847 185454
rect 393083 185218 393125 185454
rect 392805 185134 393125 185218
rect 392805 184898 392847 185134
rect 393083 184898 393125 185134
rect 392805 184866 393125 184898
rect 414874 185454 415194 185486
rect 414874 185218 414916 185454
rect 415152 185218 415194 185454
rect 414874 185134 415194 185218
rect 414874 184898 414916 185134
rect 415152 184898 415194 185134
rect 414874 184866 415194 184898
rect 420805 185454 421125 185486
rect 420805 185218 420847 185454
rect 421083 185218 421125 185454
rect 420805 185134 421125 185218
rect 420805 184898 420847 185134
rect 421083 184898 421125 185134
rect 420805 184866 421125 184898
rect 442874 185454 443194 185486
rect 442874 185218 442916 185454
rect 443152 185218 443194 185454
rect 442874 185134 443194 185218
rect 442874 184898 442916 185134
rect 443152 184898 443194 185134
rect 442874 184866 443194 184898
rect 448805 185454 449125 185486
rect 448805 185218 448847 185454
rect 449083 185218 449125 185454
rect 448805 185134 449125 185218
rect 448805 184898 448847 185134
rect 449083 184898 449125 185134
rect 448805 184866 449125 184898
rect 470874 185454 471194 185486
rect 470874 185218 470916 185454
rect 471152 185218 471194 185454
rect 470874 185134 471194 185218
rect 470874 184898 470916 185134
rect 471152 184898 471194 185134
rect 470874 184866 471194 184898
rect 476805 185454 477125 185486
rect 476805 185218 476847 185454
rect 477083 185218 477125 185454
rect 476805 185134 477125 185218
rect 476805 184898 476847 185134
rect 477083 184898 477125 185134
rect 476805 184866 477125 184898
rect 498874 185454 499194 185486
rect 498874 185218 498916 185454
rect 499152 185218 499194 185454
rect 498874 185134 499194 185218
rect 498874 184898 498916 185134
rect 499152 184898 499194 185134
rect 498874 184866 499194 184898
rect 504805 185454 505125 185486
rect 504805 185218 504847 185454
rect 505083 185218 505125 185454
rect 504805 185134 505125 185218
rect 504805 184898 504847 185134
rect 505083 184898 505125 185134
rect 504805 184866 505125 184898
rect 526874 185454 527194 185486
rect 526874 185218 526916 185454
rect 527152 185218 527194 185454
rect 526874 185134 527194 185218
rect 526874 184898 526916 185134
rect 527152 184898 527194 185134
rect 526874 184866 527194 184898
rect 532805 185454 533125 185486
rect 532805 185218 532847 185454
rect 533083 185218 533125 185454
rect 532805 185134 533125 185218
rect 532805 184898 532847 185134
rect 533083 184898 533125 185134
rect 532805 184866 533125 184898
rect 554874 185454 555194 185486
rect 554874 185218 554916 185454
rect 555152 185218 555194 185454
rect 554874 185134 555194 185218
rect 554874 184898 554916 185134
rect 555152 184898 555194 185134
rect 554874 184866 555194 184898
rect 560805 185454 561125 185486
rect 560805 185218 560847 185454
rect 561083 185218 561125 185454
rect 560805 185134 561125 185218
rect 560805 184898 560847 185134
rect 561083 184898 561125 185134
rect 560805 184866 561125 184898
rect -2006 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 -1386 161829
rect -2006 161509 -1386 161593
rect -2006 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 -1386 161509
rect -2006 134829 -1386 161273
rect 19910 161829 20230 161861
rect 19910 161593 19952 161829
rect 20188 161593 20230 161829
rect 19910 161509 20230 161593
rect 19910 161273 19952 161509
rect 20188 161273 20230 161509
rect 19910 161241 20230 161273
rect 25840 161829 26160 161861
rect 25840 161593 25882 161829
rect 26118 161593 26160 161829
rect 25840 161509 26160 161593
rect 25840 161273 25882 161509
rect 26118 161273 26160 161509
rect 25840 161241 26160 161273
rect 31771 161829 32091 161861
rect 31771 161593 31813 161829
rect 32049 161593 32091 161829
rect 31771 161509 32091 161593
rect 31771 161273 31813 161509
rect 32049 161273 32091 161509
rect 31771 161241 32091 161273
rect 47910 161829 48230 161861
rect 47910 161593 47952 161829
rect 48188 161593 48230 161829
rect 47910 161509 48230 161593
rect 47910 161273 47952 161509
rect 48188 161273 48230 161509
rect 47910 161241 48230 161273
rect 53840 161829 54160 161861
rect 53840 161593 53882 161829
rect 54118 161593 54160 161829
rect 53840 161509 54160 161593
rect 53840 161273 53882 161509
rect 54118 161273 54160 161509
rect 53840 161241 54160 161273
rect 59771 161829 60091 161861
rect 59771 161593 59813 161829
rect 60049 161593 60091 161829
rect 59771 161509 60091 161593
rect 59771 161273 59813 161509
rect 60049 161273 60091 161509
rect 59771 161241 60091 161273
rect 75910 161829 76230 161861
rect 75910 161593 75952 161829
rect 76188 161593 76230 161829
rect 75910 161509 76230 161593
rect 75910 161273 75952 161509
rect 76188 161273 76230 161509
rect 75910 161241 76230 161273
rect 81840 161829 82160 161861
rect 81840 161593 81882 161829
rect 82118 161593 82160 161829
rect 81840 161509 82160 161593
rect 81840 161273 81882 161509
rect 82118 161273 82160 161509
rect 81840 161241 82160 161273
rect 87771 161829 88091 161861
rect 87771 161593 87813 161829
rect 88049 161593 88091 161829
rect 87771 161509 88091 161593
rect 87771 161273 87813 161509
rect 88049 161273 88091 161509
rect 87771 161241 88091 161273
rect 103910 161829 104230 161861
rect 103910 161593 103952 161829
rect 104188 161593 104230 161829
rect 103910 161509 104230 161593
rect 103910 161273 103952 161509
rect 104188 161273 104230 161509
rect 103910 161241 104230 161273
rect 109840 161829 110160 161861
rect 109840 161593 109882 161829
rect 110118 161593 110160 161829
rect 109840 161509 110160 161593
rect 109840 161273 109882 161509
rect 110118 161273 110160 161509
rect 109840 161241 110160 161273
rect 115771 161829 116091 161861
rect 115771 161593 115813 161829
rect 116049 161593 116091 161829
rect 115771 161509 116091 161593
rect 115771 161273 115813 161509
rect 116049 161273 116091 161509
rect 115771 161241 116091 161273
rect 131910 161829 132230 161861
rect 131910 161593 131952 161829
rect 132188 161593 132230 161829
rect 131910 161509 132230 161593
rect 131910 161273 131952 161509
rect 132188 161273 132230 161509
rect 131910 161241 132230 161273
rect 137840 161829 138160 161861
rect 137840 161593 137882 161829
rect 138118 161593 138160 161829
rect 137840 161509 138160 161593
rect 137840 161273 137882 161509
rect 138118 161273 138160 161509
rect 137840 161241 138160 161273
rect 143771 161829 144091 161861
rect 143771 161593 143813 161829
rect 144049 161593 144091 161829
rect 143771 161509 144091 161593
rect 143771 161273 143813 161509
rect 144049 161273 144091 161509
rect 143771 161241 144091 161273
rect 159910 161829 160230 161861
rect 159910 161593 159952 161829
rect 160188 161593 160230 161829
rect 159910 161509 160230 161593
rect 159910 161273 159952 161509
rect 160188 161273 160230 161509
rect 159910 161241 160230 161273
rect 165840 161829 166160 161861
rect 165840 161593 165882 161829
rect 166118 161593 166160 161829
rect 165840 161509 166160 161593
rect 165840 161273 165882 161509
rect 166118 161273 166160 161509
rect 165840 161241 166160 161273
rect 171771 161829 172091 161861
rect 171771 161593 171813 161829
rect 172049 161593 172091 161829
rect 171771 161509 172091 161593
rect 171771 161273 171813 161509
rect 172049 161273 172091 161509
rect 171771 161241 172091 161273
rect 187910 161829 188230 161861
rect 187910 161593 187952 161829
rect 188188 161593 188230 161829
rect 187910 161509 188230 161593
rect 187910 161273 187952 161509
rect 188188 161273 188230 161509
rect 187910 161241 188230 161273
rect 193840 161829 194160 161861
rect 193840 161593 193882 161829
rect 194118 161593 194160 161829
rect 193840 161509 194160 161593
rect 193840 161273 193882 161509
rect 194118 161273 194160 161509
rect 193840 161241 194160 161273
rect 199771 161829 200091 161861
rect 199771 161593 199813 161829
rect 200049 161593 200091 161829
rect 199771 161509 200091 161593
rect 199771 161273 199813 161509
rect 200049 161273 200091 161509
rect 199771 161241 200091 161273
rect 215910 161829 216230 161861
rect 215910 161593 215952 161829
rect 216188 161593 216230 161829
rect 215910 161509 216230 161593
rect 215910 161273 215952 161509
rect 216188 161273 216230 161509
rect 215910 161241 216230 161273
rect 221840 161829 222160 161861
rect 221840 161593 221882 161829
rect 222118 161593 222160 161829
rect 221840 161509 222160 161593
rect 221840 161273 221882 161509
rect 222118 161273 222160 161509
rect 221840 161241 222160 161273
rect 227771 161829 228091 161861
rect 227771 161593 227813 161829
rect 228049 161593 228091 161829
rect 227771 161509 228091 161593
rect 227771 161273 227813 161509
rect 228049 161273 228091 161509
rect 227771 161241 228091 161273
rect 243910 161829 244230 161861
rect 243910 161593 243952 161829
rect 244188 161593 244230 161829
rect 243910 161509 244230 161593
rect 243910 161273 243952 161509
rect 244188 161273 244230 161509
rect 243910 161241 244230 161273
rect 249840 161829 250160 161861
rect 249840 161593 249882 161829
rect 250118 161593 250160 161829
rect 249840 161509 250160 161593
rect 249840 161273 249882 161509
rect 250118 161273 250160 161509
rect 249840 161241 250160 161273
rect 255771 161829 256091 161861
rect 255771 161593 255813 161829
rect 256049 161593 256091 161829
rect 255771 161509 256091 161593
rect 255771 161273 255813 161509
rect 256049 161273 256091 161509
rect 255771 161241 256091 161273
rect 271910 161829 272230 161861
rect 271910 161593 271952 161829
rect 272188 161593 272230 161829
rect 271910 161509 272230 161593
rect 271910 161273 271952 161509
rect 272188 161273 272230 161509
rect 271910 161241 272230 161273
rect 277840 161829 278160 161861
rect 277840 161593 277882 161829
rect 278118 161593 278160 161829
rect 277840 161509 278160 161593
rect 277840 161273 277882 161509
rect 278118 161273 278160 161509
rect 277840 161241 278160 161273
rect 283771 161829 284091 161861
rect 283771 161593 283813 161829
rect 284049 161593 284091 161829
rect 283771 161509 284091 161593
rect 283771 161273 283813 161509
rect 284049 161273 284091 161509
rect 283771 161241 284091 161273
rect 299910 161829 300230 161861
rect 299910 161593 299952 161829
rect 300188 161593 300230 161829
rect 299910 161509 300230 161593
rect 299910 161273 299952 161509
rect 300188 161273 300230 161509
rect 299910 161241 300230 161273
rect 305840 161829 306160 161861
rect 305840 161593 305882 161829
rect 306118 161593 306160 161829
rect 305840 161509 306160 161593
rect 305840 161273 305882 161509
rect 306118 161273 306160 161509
rect 305840 161241 306160 161273
rect 311771 161829 312091 161861
rect 311771 161593 311813 161829
rect 312049 161593 312091 161829
rect 311771 161509 312091 161593
rect 311771 161273 311813 161509
rect 312049 161273 312091 161509
rect 311771 161241 312091 161273
rect 327910 161829 328230 161861
rect 327910 161593 327952 161829
rect 328188 161593 328230 161829
rect 327910 161509 328230 161593
rect 327910 161273 327952 161509
rect 328188 161273 328230 161509
rect 327910 161241 328230 161273
rect 333840 161829 334160 161861
rect 333840 161593 333882 161829
rect 334118 161593 334160 161829
rect 333840 161509 334160 161593
rect 333840 161273 333882 161509
rect 334118 161273 334160 161509
rect 333840 161241 334160 161273
rect 339771 161829 340091 161861
rect 339771 161593 339813 161829
rect 340049 161593 340091 161829
rect 339771 161509 340091 161593
rect 339771 161273 339813 161509
rect 340049 161273 340091 161509
rect 339771 161241 340091 161273
rect 355910 161829 356230 161861
rect 355910 161593 355952 161829
rect 356188 161593 356230 161829
rect 355910 161509 356230 161593
rect 355910 161273 355952 161509
rect 356188 161273 356230 161509
rect 355910 161241 356230 161273
rect 361840 161829 362160 161861
rect 361840 161593 361882 161829
rect 362118 161593 362160 161829
rect 361840 161509 362160 161593
rect 361840 161273 361882 161509
rect 362118 161273 362160 161509
rect 361840 161241 362160 161273
rect 367771 161829 368091 161861
rect 367771 161593 367813 161829
rect 368049 161593 368091 161829
rect 367771 161509 368091 161593
rect 367771 161273 367813 161509
rect 368049 161273 368091 161509
rect 367771 161241 368091 161273
rect 383910 161829 384230 161861
rect 383910 161593 383952 161829
rect 384188 161593 384230 161829
rect 383910 161509 384230 161593
rect 383910 161273 383952 161509
rect 384188 161273 384230 161509
rect 383910 161241 384230 161273
rect 389840 161829 390160 161861
rect 389840 161593 389882 161829
rect 390118 161593 390160 161829
rect 389840 161509 390160 161593
rect 389840 161273 389882 161509
rect 390118 161273 390160 161509
rect 389840 161241 390160 161273
rect 395771 161829 396091 161861
rect 395771 161593 395813 161829
rect 396049 161593 396091 161829
rect 395771 161509 396091 161593
rect 395771 161273 395813 161509
rect 396049 161273 396091 161509
rect 395771 161241 396091 161273
rect 411910 161829 412230 161861
rect 411910 161593 411952 161829
rect 412188 161593 412230 161829
rect 411910 161509 412230 161593
rect 411910 161273 411952 161509
rect 412188 161273 412230 161509
rect 411910 161241 412230 161273
rect 417840 161829 418160 161861
rect 417840 161593 417882 161829
rect 418118 161593 418160 161829
rect 417840 161509 418160 161593
rect 417840 161273 417882 161509
rect 418118 161273 418160 161509
rect 417840 161241 418160 161273
rect 423771 161829 424091 161861
rect 423771 161593 423813 161829
rect 424049 161593 424091 161829
rect 423771 161509 424091 161593
rect 423771 161273 423813 161509
rect 424049 161273 424091 161509
rect 423771 161241 424091 161273
rect 439910 161829 440230 161861
rect 439910 161593 439952 161829
rect 440188 161593 440230 161829
rect 439910 161509 440230 161593
rect 439910 161273 439952 161509
rect 440188 161273 440230 161509
rect 439910 161241 440230 161273
rect 445840 161829 446160 161861
rect 445840 161593 445882 161829
rect 446118 161593 446160 161829
rect 445840 161509 446160 161593
rect 445840 161273 445882 161509
rect 446118 161273 446160 161509
rect 445840 161241 446160 161273
rect 451771 161829 452091 161861
rect 451771 161593 451813 161829
rect 452049 161593 452091 161829
rect 451771 161509 452091 161593
rect 451771 161273 451813 161509
rect 452049 161273 452091 161509
rect 451771 161241 452091 161273
rect 467910 161829 468230 161861
rect 467910 161593 467952 161829
rect 468188 161593 468230 161829
rect 467910 161509 468230 161593
rect 467910 161273 467952 161509
rect 468188 161273 468230 161509
rect 467910 161241 468230 161273
rect 473840 161829 474160 161861
rect 473840 161593 473882 161829
rect 474118 161593 474160 161829
rect 473840 161509 474160 161593
rect 473840 161273 473882 161509
rect 474118 161273 474160 161509
rect 473840 161241 474160 161273
rect 479771 161829 480091 161861
rect 479771 161593 479813 161829
rect 480049 161593 480091 161829
rect 479771 161509 480091 161593
rect 479771 161273 479813 161509
rect 480049 161273 480091 161509
rect 479771 161241 480091 161273
rect 495910 161829 496230 161861
rect 495910 161593 495952 161829
rect 496188 161593 496230 161829
rect 495910 161509 496230 161593
rect 495910 161273 495952 161509
rect 496188 161273 496230 161509
rect 495910 161241 496230 161273
rect 501840 161829 502160 161861
rect 501840 161593 501882 161829
rect 502118 161593 502160 161829
rect 501840 161509 502160 161593
rect 501840 161273 501882 161509
rect 502118 161273 502160 161509
rect 501840 161241 502160 161273
rect 507771 161829 508091 161861
rect 507771 161593 507813 161829
rect 508049 161593 508091 161829
rect 507771 161509 508091 161593
rect 507771 161273 507813 161509
rect 508049 161273 508091 161509
rect 507771 161241 508091 161273
rect 523910 161829 524230 161861
rect 523910 161593 523952 161829
rect 524188 161593 524230 161829
rect 523910 161509 524230 161593
rect 523910 161273 523952 161509
rect 524188 161273 524230 161509
rect 523910 161241 524230 161273
rect 529840 161829 530160 161861
rect 529840 161593 529882 161829
rect 530118 161593 530160 161829
rect 529840 161509 530160 161593
rect 529840 161273 529882 161509
rect 530118 161273 530160 161509
rect 529840 161241 530160 161273
rect 535771 161829 536091 161861
rect 535771 161593 535813 161829
rect 536049 161593 536091 161829
rect 535771 161509 536091 161593
rect 535771 161273 535813 161509
rect 536049 161273 536091 161509
rect 535771 161241 536091 161273
rect 551910 161829 552230 161861
rect 551910 161593 551952 161829
rect 552188 161593 552230 161829
rect 551910 161509 552230 161593
rect 551910 161273 551952 161509
rect 552188 161273 552230 161509
rect 551910 161241 552230 161273
rect 557840 161829 558160 161861
rect 557840 161593 557882 161829
rect 558118 161593 558160 161829
rect 557840 161509 558160 161593
rect 557840 161273 557882 161509
rect 558118 161273 558160 161509
rect 557840 161241 558160 161273
rect 563771 161829 564091 161861
rect 563771 161593 563813 161829
rect 564049 161593 564091 161829
rect 563771 161509 564091 161593
rect 563771 161273 563813 161509
rect 564049 161273 564091 161509
rect 563771 161241 564091 161273
rect 573494 161829 574114 188273
rect 573494 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 574114 161829
rect 573494 161509 574114 161593
rect 573494 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 574114 161509
rect 22874 158454 23194 158486
rect 22874 158218 22916 158454
rect 23152 158218 23194 158454
rect 22874 158134 23194 158218
rect 22874 157898 22916 158134
rect 23152 157898 23194 158134
rect 22874 157866 23194 157898
rect 28805 158454 29125 158486
rect 28805 158218 28847 158454
rect 29083 158218 29125 158454
rect 28805 158134 29125 158218
rect 28805 157898 28847 158134
rect 29083 157898 29125 158134
rect 28805 157866 29125 157898
rect 50874 158454 51194 158486
rect 50874 158218 50916 158454
rect 51152 158218 51194 158454
rect 50874 158134 51194 158218
rect 50874 157898 50916 158134
rect 51152 157898 51194 158134
rect 50874 157866 51194 157898
rect 56805 158454 57125 158486
rect 56805 158218 56847 158454
rect 57083 158218 57125 158454
rect 56805 158134 57125 158218
rect 56805 157898 56847 158134
rect 57083 157898 57125 158134
rect 56805 157866 57125 157898
rect 78874 158454 79194 158486
rect 78874 158218 78916 158454
rect 79152 158218 79194 158454
rect 78874 158134 79194 158218
rect 78874 157898 78916 158134
rect 79152 157898 79194 158134
rect 78874 157866 79194 157898
rect 84805 158454 85125 158486
rect 84805 158218 84847 158454
rect 85083 158218 85125 158454
rect 84805 158134 85125 158218
rect 84805 157898 84847 158134
rect 85083 157898 85125 158134
rect 84805 157866 85125 157898
rect 106874 158454 107194 158486
rect 106874 158218 106916 158454
rect 107152 158218 107194 158454
rect 106874 158134 107194 158218
rect 106874 157898 106916 158134
rect 107152 157898 107194 158134
rect 106874 157866 107194 157898
rect 112805 158454 113125 158486
rect 112805 158218 112847 158454
rect 113083 158218 113125 158454
rect 112805 158134 113125 158218
rect 112805 157898 112847 158134
rect 113083 157898 113125 158134
rect 112805 157866 113125 157898
rect 134874 158454 135194 158486
rect 134874 158218 134916 158454
rect 135152 158218 135194 158454
rect 134874 158134 135194 158218
rect 134874 157898 134916 158134
rect 135152 157898 135194 158134
rect 134874 157866 135194 157898
rect 140805 158454 141125 158486
rect 140805 158218 140847 158454
rect 141083 158218 141125 158454
rect 140805 158134 141125 158218
rect 140805 157898 140847 158134
rect 141083 157898 141125 158134
rect 140805 157866 141125 157898
rect 162874 158454 163194 158486
rect 162874 158218 162916 158454
rect 163152 158218 163194 158454
rect 162874 158134 163194 158218
rect 162874 157898 162916 158134
rect 163152 157898 163194 158134
rect 162874 157866 163194 157898
rect 168805 158454 169125 158486
rect 168805 158218 168847 158454
rect 169083 158218 169125 158454
rect 168805 158134 169125 158218
rect 168805 157898 168847 158134
rect 169083 157898 169125 158134
rect 168805 157866 169125 157898
rect 190874 158454 191194 158486
rect 190874 158218 190916 158454
rect 191152 158218 191194 158454
rect 190874 158134 191194 158218
rect 190874 157898 190916 158134
rect 191152 157898 191194 158134
rect 190874 157866 191194 157898
rect 196805 158454 197125 158486
rect 196805 158218 196847 158454
rect 197083 158218 197125 158454
rect 196805 158134 197125 158218
rect 196805 157898 196847 158134
rect 197083 157898 197125 158134
rect 196805 157866 197125 157898
rect 218874 158454 219194 158486
rect 218874 158218 218916 158454
rect 219152 158218 219194 158454
rect 218874 158134 219194 158218
rect 218874 157898 218916 158134
rect 219152 157898 219194 158134
rect 218874 157866 219194 157898
rect 224805 158454 225125 158486
rect 224805 158218 224847 158454
rect 225083 158218 225125 158454
rect 224805 158134 225125 158218
rect 224805 157898 224847 158134
rect 225083 157898 225125 158134
rect 224805 157866 225125 157898
rect 246874 158454 247194 158486
rect 246874 158218 246916 158454
rect 247152 158218 247194 158454
rect 246874 158134 247194 158218
rect 246874 157898 246916 158134
rect 247152 157898 247194 158134
rect 246874 157866 247194 157898
rect 252805 158454 253125 158486
rect 252805 158218 252847 158454
rect 253083 158218 253125 158454
rect 252805 158134 253125 158218
rect 252805 157898 252847 158134
rect 253083 157898 253125 158134
rect 252805 157866 253125 157898
rect 274874 158454 275194 158486
rect 274874 158218 274916 158454
rect 275152 158218 275194 158454
rect 274874 158134 275194 158218
rect 274874 157898 274916 158134
rect 275152 157898 275194 158134
rect 274874 157866 275194 157898
rect 280805 158454 281125 158486
rect 280805 158218 280847 158454
rect 281083 158218 281125 158454
rect 280805 158134 281125 158218
rect 280805 157898 280847 158134
rect 281083 157898 281125 158134
rect 280805 157866 281125 157898
rect 302874 158454 303194 158486
rect 302874 158218 302916 158454
rect 303152 158218 303194 158454
rect 302874 158134 303194 158218
rect 302874 157898 302916 158134
rect 303152 157898 303194 158134
rect 302874 157866 303194 157898
rect 308805 158454 309125 158486
rect 308805 158218 308847 158454
rect 309083 158218 309125 158454
rect 308805 158134 309125 158218
rect 308805 157898 308847 158134
rect 309083 157898 309125 158134
rect 308805 157866 309125 157898
rect 330874 158454 331194 158486
rect 330874 158218 330916 158454
rect 331152 158218 331194 158454
rect 330874 158134 331194 158218
rect 330874 157898 330916 158134
rect 331152 157898 331194 158134
rect 330874 157866 331194 157898
rect 336805 158454 337125 158486
rect 336805 158218 336847 158454
rect 337083 158218 337125 158454
rect 336805 158134 337125 158218
rect 336805 157898 336847 158134
rect 337083 157898 337125 158134
rect 336805 157866 337125 157898
rect 358874 158454 359194 158486
rect 358874 158218 358916 158454
rect 359152 158218 359194 158454
rect 358874 158134 359194 158218
rect 358874 157898 358916 158134
rect 359152 157898 359194 158134
rect 358874 157866 359194 157898
rect 364805 158454 365125 158486
rect 364805 158218 364847 158454
rect 365083 158218 365125 158454
rect 364805 158134 365125 158218
rect 364805 157898 364847 158134
rect 365083 157898 365125 158134
rect 364805 157866 365125 157898
rect 386874 158454 387194 158486
rect 386874 158218 386916 158454
rect 387152 158218 387194 158454
rect 386874 158134 387194 158218
rect 386874 157898 386916 158134
rect 387152 157898 387194 158134
rect 386874 157866 387194 157898
rect 392805 158454 393125 158486
rect 392805 158218 392847 158454
rect 393083 158218 393125 158454
rect 392805 158134 393125 158218
rect 392805 157898 392847 158134
rect 393083 157898 393125 158134
rect 392805 157866 393125 157898
rect 414874 158454 415194 158486
rect 414874 158218 414916 158454
rect 415152 158218 415194 158454
rect 414874 158134 415194 158218
rect 414874 157898 414916 158134
rect 415152 157898 415194 158134
rect 414874 157866 415194 157898
rect 420805 158454 421125 158486
rect 420805 158218 420847 158454
rect 421083 158218 421125 158454
rect 420805 158134 421125 158218
rect 420805 157898 420847 158134
rect 421083 157898 421125 158134
rect 420805 157866 421125 157898
rect 442874 158454 443194 158486
rect 442874 158218 442916 158454
rect 443152 158218 443194 158454
rect 442874 158134 443194 158218
rect 442874 157898 442916 158134
rect 443152 157898 443194 158134
rect 442874 157866 443194 157898
rect 448805 158454 449125 158486
rect 448805 158218 448847 158454
rect 449083 158218 449125 158454
rect 448805 158134 449125 158218
rect 448805 157898 448847 158134
rect 449083 157898 449125 158134
rect 448805 157866 449125 157898
rect 470874 158454 471194 158486
rect 470874 158218 470916 158454
rect 471152 158218 471194 158454
rect 470874 158134 471194 158218
rect 470874 157898 470916 158134
rect 471152 157898 471194 158134
rect 470874 157866 471194 157898
rect 476805 158454 477125 158486
rect 476805 158218 476847 158454
rect 477083 158218 477125 158454
rect 476805 158134 477125 158218
rect 476805 157898 476847 158134
rect 477083 157898 477125 158134
rect 476805 157866 477125 157898
rect 498874 158454 499194 158486
rect 498874 158218 498916 158454
rect 499152 158218 499194 158454
rect 498874 158134 499194 158218
rect 498874 157898 498916 158134
rect 499152 157898 499194 158134
rect 498874 157866 499194 157898
rect 504805 158454 505125 158486
rect 504805 158218 504847 158454
rect 505083 158218 505125 158454
rect 504805 158134 505125 158218
rect 504805 157898 504847 158134
rect 505083 157898 505125 158134
rect 504805 157866 505125 157898
rect 526874 158454 527194 158486
rect 526874 158218 526916 158454
rect 527152 158218 527194 158454
rect 526874 158134 527194 158218
rect 526874 157898 526916 158134
rect 527152 157898 527194 158134
rect 526874 157866 527194 157898
rect 532805 158454 533125 158486
rect 532805 158218 532847 158454
rect 533083 158218 533125 158454
rect 532805 158134 533125 158218
rect 532805 157898 532847 158134
rect 533083 157898 533125 158134
rect 532805 157866 533125 157898
rect 554874 158454 555194 158486
rect 554874 158218 554916 158454
rect 555152 158218 555194 158454
rect 554874 158134 555194 158218
rect 554874 157898 554916 158134
rect 555152 157898 555194 158134
rect 554874 157866 555194 157898
rect 560805 158454 561125 158486
rect 560805 158218 560847 158454
rect 561083 158218 561125 158454
rect 560805 158134 561125 158218
rect 560805 157898 560847 158134
rect 561083 157898 561125 158134
rect 560805 157866 561125 157898
rect -2006 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 -1386 134829
rect -2006 134509 -1386 134593
rect -2006 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 -1386 134509
rect -2006 107829 -1386 134273
rect 19910 134829 20230 134861
rect 19910 134593 19952 134829
rect 20188 134593 20230 134829
rect 19910 134509 20230 134593
rect 19910 134273 19952 134509
rect 20188 134273 20230 134509
rect 19910 134241 20230 134273
rect 25840 134829 26160 134861
rect 25840 134593 25882 134829
rect 26118 134593 26160 134829
rect 25840 134509 26160 134593
rect 25840 134273 25882 134509
rect 26118 134273 26160 134509
rect 25840 134241 26160 134273
rect 31771 134829 32091 134861
rect 31771 134593 31813 134829
rect 32049 134593 32091 134829
rect 31771 134509 32091 134593
rect 31771 134273 31813 134509
rect 32049 134273 32091 134509
rect 31771 134241 32091 134273
rect 47910 134829 48230 134861
rect 47910 134593 47952 134829
rect 48188 134593 48230 134829
rect 47910 134509 48230 134593
rect 47910 134273 47952 134509
rect 48188 134273 48230 134509
rect 47910 134241 48230 134273
rect 53840 134829 54160 134861
rect 53840 134593 53882 134829
rect 54118 134593 54160 134829
rect 53840 134509 54160 134593
rect 53840 134273 53882 134509
rect 54118 134273 54160 134509
rect 53840 134241 54160 134273
rect 59771 134829 60091 134861
rect 59771 134593 59813 134829
rect 60049 134593 60091 134829
rect 59771 134509 60091 134593
rect 59771 134273 59813 134509
rect 60049 134273 60091 134509
rect 59771 134241 60091 134273
rect 75910 134829 76230 134861
rect 75910 134593 75952 134829
rect 76188 134593 76230 134829
rect 75910 134509 76230 134593
rect 75910 134273 75952 134509
rect 76188 134273 76230 134509
rect 75910 134241 76230 134273
rect 81840 134829 82160 134861
rect 81840 134593 81882 134829
rect 82118 134593 82160 134829
rect 81840 134509 82160 134593
rect 81840 134273 81882 134509
rect 82118 134273 82160 134509
rect 81840 134241 82160 134273
rect 87771 134829 88091 134861
rect 87771 134593 87813 134829
rect 88049 134593 88091 134829
rect 87771 134509 88091 134593
rect 87771 134273 87813 134509
rect 88049 134273 88091 134509
rect 87771 134241 88091 134273
rect 103910 134829 104230 134861
rect 103910 134593 103952 134829
rect 104188 134593 104230 134829
rect 103910 134509 104230 134593
rect 103910 134273 103952 134509
rect 104188 134273 104230 134509
rect 103910 134241 104230 134273
rect 109840 134829 110160 134861
rect 109840 134593 109882 134829
rect 110118 134593 110160 134829
rect 109840 134509 110160 134593
rect 109840 134273 109882 134509
rect 110118 134273 110160 134509
rect 109840 134241 110160 134273
rect 115771 134829 116091 134861
rect 115771 134593 115813 134829
rect 116049 134593 116091 134829
rect 115771 134509 116091 134593
rect 115771 134273 115813 134509
rect 116049 134273 116091 134509
rect 115771 134241 116091 134273
rect 131910 134829 132230 134861
rect 131910 134593 131952 134829
rect 132188 134593 132230 134829
rect 131910 134509 132230 134593
rect 131910 134273 131952 134509
rect 132188 134273 132230 134509
rect 131910 134241 132230 134273
rect 137840 134829 138160 134861
rect 137840 134593 137882 134829
rect 138118 134593 138160 134829
rect 137840 134509 138160 134593
rect 137840 134273 137882 134509
rect 138118 134273 138160 134509
rect 137840 134241 138160 134273
rect 143771 134829 144091 134861
rect 143771 134593 143813 134829
rect 144049 134593 144091 134829
rect 143771 134509 144091 134593
rect 143771 134273 143813 134509
rect 144049 134273 144091 134509
rect 143771 134241 144091 134273
rect 159910 134829 160230 134861
rect 159910 134593 159952 134829
rect 160188 134593 160230 134829
rect 159910 134509 160230 134593
rect 159910 134273 159952 134509
rect 160188 134273 160230 134509
rect 159910 134241 160230 134273
rect 165840 134829 166160 134861
rect 165840 134593 165882 134829
rect 166118 134593 166160 134829
rect 165840 134509 166160 134593
rect 165840 134273 165882 134509
rect 166118 134273 166160 134509
rect 165840 134241 166160 134273
rect 171771 134829 172091 134861
rect 171771 134593 171813 134829
rect 172049 134593 172091 134829
rect 171771 134509 172091 134593
rect 171771 134273 171813 134509
rect 172049 134273 172091 134509
rect 171771 134241 172091 134273
rect 187910 134829 188230 134861
rect 187910 134593 187952 134829
rect 188188 134593 188230 134829
rect 187910 134509 188230 134593
rect 187910 134273 187952 134509
rect 188188 134273 188230 134509
rect 187910 134241 188230 134273
rect 193840 134829 194160 134861
rect 193840 134593 193882 134829
rect 194118 134593 194160 134829
rect 193840 134509 194160 134593
rect 193840 134273 193882 134509
rect 194118 134273 194160 134509
rect 193840 134241 194160 134273
rect 199771 134829 200091 134861
rect 199771 134593 199813 134829
rect 200049 134593 200091 134829
rect 199771 134509 200091 134593
rect 199771 134273 199813 134509
rect 200049 134273 200091 134509
rect 199771 134241 200091 134273
rect 215910 134829 216230 134861
rect 215910 134593 215952 134829
rect 216188 134593 216230 134829
rect 215910 134509 216230 134593
rect 215910 134273 215952 134509
rect 216188 134273 216230 134509
rect 215910 134241 216230 134273
rect 221840 134829 222160 134861
rect 221840 134593 221882 134829
rect 222118 134593 222160 134829
rect 221840 134509 222160 134593
rect 221840 134273 221882 134509
rect 222118 134273 222160 134509
rect 221840 134241 222160 134273
rect 227771 134829 228091 134861
rect 227771 134593 227813 134829
rect 228049 134593 228091 134829
rect 227771 134509 228091 134593
rect 227771 134273 227813 134509
rect 228049 134273 228091 134509
rect 227771 134241 228091 134273
rect 243910 134829 244230 134861
rect 243910 134593 243952 134829
rect 244188 134593 244230 134829
rect 243910 134509 244230 134593
rect 243910 134273 243952 134509
rect 244188 134273 244230 134509
rect 243910 134241 244230 134273
rect 249840 134829 250160 134861
rect 249840 134593 249882 134829
rect 250118 134593 250160 134829
rect 249840 134509 250160 134593
rect 249840 134273 249882 134509
rect 250118 134273 250160 134509
rect 249840 134241 250160 134273
rect 255771 134829 256091 134861
rect 255771 134593 255813 134829
rect 256049 134593 256091 134829
rect 255771 134509 256091 134593
rect 255771 134273 255813 134509
rect 256049 134273 256091 134509
rect 255771 134241 256091 134273
rect 271910 134829 272230 134861
rect 271910 134593 271952 134829
rect 272188 134593 272230 134829
rect 271910 134509 272230 134593
rect 271910 134273 271952 134509
rect 272188 134273 272230 134509
rect 271910 134241 272230 134273
rect 277840 134829 278160 134861
rect 277840 134593 277882 134829
rect 278118 134593 278160 134829
rect 277840 134509 278160 134593
rect 277840 134273 277882 134509
rect 278118 134273 278160 134509
rect 277840 134241 278160 134273
rect 283771 134829 284091 134861
rect 283771 134593 283813 134829
rect 284049 134593 284091 134829
rect 283771 134509 284091 134593
rect 283771 134273 283813 134509
rect 284049 134273 284091 134509
rect 283771 134241 284091 134273
rect 299910 134829 300230 134861
rect 299910 134593 299952 134829
rect 300188 134593 300230 134829
rect 299910 134509 300230 134593
rect 299910 134273 299952 134509
rect 300188 134273 300230 134509
rect 299910 134241 300230 134273
rect 305840 134829 306160 134861
rect 305840 134593 305882 134829
rect 306118 134593 306160 134829
rect 305840 134509 306160 134593
rect 305840 134273 305882 134509
rect 306118 134273 306160 134509
rect 305840 134241 306160 134273
rect 311771 134829 312091 134861
rect 311771 134593 311813 134829
rect 312049 134593 312091 134829
rect 311771 134509 312091 134593
rect 311771 134273 311813 134509
rect 312049 134273 312091 134509
rect 311771 134241 312091 134273
rect 327910 134829 328230 134861
rect 327910 134593 327952 134829
rect 328188 134593 328230 134829
rect 327910 134509 328230 134593
rect 327910 134273 327952 134509
rect 328188 134273 328230 134509
rect 327910 134241 328230 134273
rect 333840 134829 334160 134861
rect 333840 134593 333882 134829
rect 334118 134593 334160 134829
rect 333840 134509 334160 134593
rect 333840 134273 333882 134509
rect 334118 134273 334160 134509
rect 333840 134241 334160 134273
rect 339771 134829 340091 134861
rect 339771 134593 339813 134829
rect 340049 134593 340091 134829
rect 339771 134509 340091 134593
rect 339771 134273 339813 134509
rect 340049 134273 340091 134509
rect 339771 134241 340091 134273
rect 355910 134829 356230 134861
rect 355910 134593 355952 134829
rect 356188 134593 356230 134829
rect 355910 134509 356230 134593
rect 355910 134273 355952 134509
rect 356188 134273 356230 134509
rect 355910 134241 356230 134273
rect 361840 134829 362160 134861
rect 361840 134593 361882 134829
rect 362118 134593 362160 134829
rect 361840 134509 362160 134593
rect 361840 134273 361882 134509
rect 362118 134273 362160 134509
rect 361840 134241 362160 134273
rect 367771 134829 368091 134861
rect 367771 134593 367813 134829
rect 368049 134593 368091 134829
rect 367771 134509 368091 134593
rect 367771 134273 367813 134509
rect 368049 134273 368091 134509
rect 367771 134241 368091 134273
rect 383910 134829 384230 134861
rect 383910 134593 383952 134829
rect 384188 134593 384230 134829
rect 383910 134509 384230 134593
rect 383910 134273 383952 134509
rect 384188 134273 384230 134509
rect 383910 134241 384230 134273
rect 389840 134829 390160 134861
rect 389840 134593 389882 134829
rect 390118 134593 390160 134829
rect 389840 134509 390160 134593
rect 389840 134273 389882 134509
rect 390118 134273 390160 134509
rect 389840 134241 390160 134273
rect 395771 134829 396091 134861
rect 395771 134593 395813 134829
rect 396049 134593 396091 134829
rect 395771 134509 396091 134593
rect 395771 134273 395813 134509
rect 396049 134273 396091 134509
rect 395771 134241 396091 134273
rect 411910 134829 412230 134861
rect 411910 134593 411952 134829
rect 412188 134593 412230 134829
rect 411910 134509 412230 134593
rect 411910 134273 411952 134509
rect 412188 134273 412230 134509
rect 411910 134241 412230 134273
rect 417840 134829 418160 134861
rect 417840 134593 417882 134829
rect 418118 134593 418160 134829
rect 417840 134509 418160 134593
rect 417840 134273 417882 134509
rect 418118 134273 418160 134509
rect 417840 134241 418160 134273
rect 423771 134829 424091 134861
rect 423771 134593 423813 134829
rect 424049 134593 424091 134829
rect 423771 134509 424091 134593
rect 423771 134273 423813 134509
rect 424049 134273 424091 134509
rect 423771 134241 424091 134273
rect 439910 134829 440230 134861
rect 439910 134593 439952 134829
rect 440188 134593 440230 134829
rect 439910 134509 440230 134593
rect 439910 134273 439952 134509
rect 440188 134273 440230 134509
rect 439910 134241 440230 134273
rect 445840 134829 446160 134861
rect 445840 134593 445882 134829
rect 446118 134593 446160 134829
rect 445840 134509 446160 134593
rect 445840 134273 445882 134509
rect 446118 134273 446160 134509
rect 445840 134241 446160 134273
rect 451771 134829 452091 134861
rect 451771 134593 451813 134829
rect 452049 134593 452091 134829
rect 451771 134509 452091 134593
rect 451771 134273 451813 134509
rect 452049 134273 452091 134509
rect 451771 134241 452091 134273
rect 467910 134829 468230 134861
rect 467910 134593 467952 134829
rect 468188 134593 468230 134829
rect 467910 134509 468230 134593
rect 467910 134273 467952 134509
rect 468188 134273 468230 134509
rect 467910 134241 468230 134273
rect 473840 134829 474160 134861
rect 473840 134593 473882 134829
rect 474118 134593 474160 134829
rect 473840 134509 474160 134593
rect 473840 134273 473882 134509
rect 474118 134273 474160 134509
rect 473840 134241 474160 134273
rect 479771 134829 480091 134861
rect 479771 134593 479813 134829
rect 480049 134593 480091 134829
rect 479771 134509 480091 134593
rect 479771 134273 479813 134509
rect 480049 134273 480091 134509
rect 479771 134241 480091 134273
rect 495910 134829 496230 134861
rect 495910 134593 495952 134829
rect 496188 134593 496230 134829
rect 495910 134509 496230 134593
rect 495910 134273 495952 134509
rect 496188 134273 496230 134509
rect 495910 134241 496230 134273
rect 501840 134829 502160 134861
rect 501840 134593 501882 134829
rect 502118 134593 502160 134829
rect 501840 134509 502160 134593
rect 501840 134273 501882 134509
rect 502118 134273 502160 134509
rect 501840 134241 502160 134273
rect 507771 134829 508091 134861
rect 507771 134593 507813 134829
rect 508049 134593 508091 134829
rect 507771 134509 508091 134593
rect 507771 134273 507813 134509
rect 508049 134273 508091 134509
rect 507771 134241 508091 134273
rect 523910 134829 524230 134861
rect 523910 134593 523952 134829
rect 524188 134593 524230 134829
rect 523910 134509 524230 134593
rect 523910 134273 523952 134509
rect 524188 134273 524230 134509
rect 523910 134241 524230 134273
rect 529840 134829 530160 134861
rect 529840 134593 529882 134829
rect 530118 134593 530160 134829
rect 529840 134509 530160 134593
rect 529840 134273 529882 134509
rect 530118 134273 530160 134509
rect 529840 134241 530160 134273
rect 535771 134829 536091 134861
rect 535771 134593 535813 134829
rect 536049 134593 536091 134829
rect 535771 134509 536091 134593
rect 535771 134273 535813 134509
rect 536049 134273 536091 134509
rect 535771 134241 536091 134273
rect 551910 134829 552230 134861
rect 551910 134593 551952 134829
rect 552188 134593 552230 134829
rect 551910 134509 552230 134593
rect 551910 134273 551952 134509
rect 552188 134273 552230 134509
rect 551910 134241 552230 134273
rect 557840 134829 558160 134861
rect 557840 134593 557882 134829
rect 558118 134593 558160 134829
rect 557840 134509 558160 134593
rect 557840 134273 557882 134509
rect 558118 134273 558160 134509
rect 557840 134241 558160 134273
rect 563771 134829 564091 134861
rect 563771 134593 563813 134829
rect 564049 134593 564091 134829
rect 563771 134509 564091 134593
rect 563771 134273 563813 134509
rect 564049 134273 564091 134509
rect 563771 134241 564091 134273
rect 573494 134829 574114 161273
rect 573494 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 574114 134829
rect 573494 134509 574114 134593
rect 573494 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 574114 134509
rect 22874 131454 23194 131486
rect 22874 131218 22916 131454
rect 23152 131218 23194 131454
rect 22874 131134 23194 131218
rect 22874 130898 22916 131134
rect 23152 130898 23194 131134
rect 22874 130866 23194 130898
rect 28805 131454 29125 131486
rect 28805 131218 28847 131454
rect 29083 131218 29125 131454
rect 28805 131134 29125 131218
rect 28805 130898 28847 131134
rect 29083 130898 29125 131134
rect 28805 130866 29125 130898
rect 50874 131454 51194 131486
rect 50874 131218 50916 131454
rect 51152 131218 51194 131454
rect 50874 131134 51194 131218
rect 50874 130898 50916 131134
rect 51152 130898 51194 131134
rect 50874 130866 51194 130898
rect 56805 131454 57125 131486
rect 56805 131218 56847 131454
rect 57083 131218 57125 131454
rect 56805 131134 57125 131218
rect 56805 130898 56847 131134
rect 57083 130898 57125 131134
rect 56805 130866 57125 130898
rect 78874 131454 79194 131486
rect 78874 131218 78916 131454
rect 79152 131218 79194 131454
rect 78874 131134 79194 131218
rect 78874 130898 78916 131134
rect 79152 130898 79194 131134
rect 78874 130866 79194 130898
rect 84805 131454 85125 131486
rect 84805 131218 84847 131454
rect 85083 131218 85125 131454
rect 84805 131134 85125 131218
rect 84805 130898 84847 131134
rect 85083 130898 85125 131134
rect 84805 130866 85125 130898
rect 106874 131454 107194 131486
rect 106874 131218 106916 131454
rect 107152 131218 107194 131454
rect 106874 131134 107194 131218
rect 106874 130898 106916 131134
rect 107152 130898 107194 131134
rect 106874 130866 107194 130898
rect 112805 131454 113125 131486
rect 112805 131218 112847 131454
rect 113083 131218 113125 131454
rect 112805 131134 113125 131218
rect 112805 130898 112847 131134
rect 113083 130898 113125 131134
rect 112805 130866 113125 130898
rect 134874 131454 135194 131486
rect 134874 131218 134916 131454
rect 135152 131218 135194 131454
rect 134874 131134 135194 131218
rect 134874 130898 134916 131134
rect 135152 130898 135194 131134
rect 134874 130866 135194 130898
rect 140805 131454 141125 131486
rect 140805 131218 140847 131454
rect 141083 131218 141125 131454
rect 140805 131134 141125 131218
rect 140805 130898 140847 131134
rect 141083 130898 141125 131134
rect 140805 130866 141125 130898
rect 162874 131454 163194 131486
rect 162874 131218 162916 131454
rect 163152 131218 163194 131454
rect 162874 131134 163194 131218
rect 162874 130898 162916 131134
rect 163152 130898 163194 131134
rect 162874 130866 163194 130898
rect 168805 131454 169125 131486
rect 168805 131218 168847 131454
rect 169083 131218 169125 131454
rect 168805 131134 169125 131218
rect 168805 130898 168847 131134
rect 169083 130898 169125 131134
rect 168805 130866 169125 130898
rect 190874 131454 191194 131486
rect 190874 131218 190916 131454
rect 191152 131218 191194 131454
rect 190874 131134 191194 131218
rect 190874 130898 190916 131134
rect 191152 130898 191194 131134
rect 190874 130866 191194 130898
rect 196805 131454 197125 131486
rect 196805 131218 196847 131454
rect 197083 131218 197125 131454
rect 196805 131134 197125 131218
rect 196805 130898 196847 131134
rect 197083 130898 197125 131134
rect 196805 130866 197125 130898
rect 218874 131454 219194 131486
rect 218874 131218 218916 131454
rect 219152 131218 219194 131454
rect 218874 131134 219194 131218
rect 218874 130898 218916 131134
rect 219152 130898 219194 131134
rect 218874 130866 219194 130898
rect 224805 131454 225125 131486
rect 224805 131218 224847 131454
rect 225083 131218 225125 131454
rect 224805 131134 225125 131218
rect 224805 130898 224847 131134
rect 225083 130898 225125 131134
rect 224805 130866 225125 130898
rect 246874 131454 247194 131486
rect 246874 131218 246916 131454
rect 247152 131218 247194 131454
rect 246874 131134 247194 131218
rect 246874 130898 246916 131134
rect 247152 130898 247194 131134
rect 246874 130866 247194 130898
rect 252805 131454 253125 131486
rect 252805 131218 252847 131454
rect 253083 131218 253125 131454
rect 252805 131134 253125 131218
rect 252805 130898 252847 131134
rect 253083 130898 253125 131134
rect 252805 130866 253125 130898
rect 274874 131454 275194 131486
rect 274874 131218 274916 131454
rect 275152 131218 275194 131454
rect 274874 131134 275194 131218
rect 274874 130898 274916 131134
rect 275152 130898 275194 131134
rect 274874 130866 275194 130898
rect 280805 131454 281125 131486
rect 280805 131218 280847 131454
rect 281083 131218 281125 131454
rect 280805 131134 281125 131218
rect 280805 130898 280847 131134
rect 281083 130898 281125 131134
rect 280805 130866 281125 130898
rect 302874 131454 303194 131486
rect 302874 131218 302916 131454
rect 303152 131218 303194 131454
rect 302874 131134 303194 131218
rect 302874 130898 302916 131134
rect 303152 130898 303194 131134
rect 302874 130866 303194 130898
rect 308805 131454 309125 131486
rect 308805 131218 308847 131454
rect 309083 131218 309125 131454
rect 308805 131134 309125 131218
rect 308805 130898 308847 131134
rect 309083 130898 309125 131134
rect 308805 130866 309125 130898
rect 330874 131454 331194 131486
rect 330874 131218 330916 131454
rect 331152 131218 331194 131454
rect 330874 131134 331194 131218
rect 330874 130898 330916 131134
rect 331152 130898 331194 131134
rect 330874 130866 331194 130898
rect 336805 131454 337125 131486
rect 336805 131218 336847 131454
rect 337083 131218 337125 131454
rect 336805 131134 337125 131218
rect 336805 130898 336847 131134
rect 337083 130898 337125 131134
rect 336805 130866 337125 130898
rect 358874 131454 359194 131486
rect 358874 131218 358916 131454
rect 359152 131218 359194 131454
rect 358874 131134 359194 131218
rect 358874 130898 358916 131134
rect 359152 130898 359194 131134
rect 358874 130866 359194 130898
rect 364805 131454 365125 131486
rect 364805 131218 364847 131454
rect 365083 131218 365125 131454
rect 364805 131134 365125 131218
rect 364805 130898 364847 131134
rect 365083 130898 365125 131134
rect 364805 130866 365125 130898
rect 386874 131454 387194 131486
rect 386874 131218 386916 131454
rect 387152 131218 387194 131454
rect 386874 131134 387194 131218
rect 386874 130898 386916 131134
rect 387152 130898 387194 131134
rect 386874 130866 387194 130898
rect 392805 131454 393125 131486
rect 392805 131218 392847 131454
rect 393083 131218 393125 131454
rect 392805 131134 393125 131218
rect 392805 130898 392847 131134
rect 393083 130898 393125 131134
rect 392805 130866 393125 130898
rect 414874 131454 415194 131486
rect 414874 131218 414916 131454
rect 415152 131218 415194 131454
rect 414874 131134 415194 131218
rect 414874 130898 414916 131134
rect 415152 130898 415194 131134
rect 414874 130866 415194 130898
rect 420805 131454 421125 131486
rect 420805 131218 420847 131454
rect 421083 131218 421125 131454
rect 420805 131134 421125 131218
rect 420805 130898 420847 131134
rect 421083 130898 421125 131134
rect 420805 130866 421125 130898
rect 442874 131454 443194 131486
rect 442874 131218 442916 131454
rect 443152 131218 443194 131454
rect 442874 131134 443194 131218
rect 442874 130898 442916 131134
rect 443152 130898 443194 131134
rect 442874 130866 443194 130898
rect 448805 131454 449125 131486
rect 448805 131218 448847 131454
rect 449083 131218 449125 131454
rect 448805 131134 449125 131218
rect 448805 130898 448847 131134
rect 449083 130898 449125 131134
rect 448805 130866 449125 130898
rect 470874 131454 471194 131486
rect 470874 131218 470916 131454
rect 471152 131218 471194 131454
rect 470874 131134 471194 131218
rect 470874 130898 470916 131134
rect 471152 130898 471194 131134
rect 470874 130866 471194 130898
rect 476805 131454 477125 131486
rect 476805 131218 476847 131454
rect 477083 131218 477125 131454
rect 476805 131134 477125 131218
rect 476805 130898 476847 131134
rect 477083 130898 477125 131134
rect 476805 130866 477125 130898
rect 498874 131454 499194 131486
rect 498874 131218 498916 131454
rect 499152 131218 499194 131454
rect 498874 131134 499194 131218
rect 498874 130898 498916 131134
rect 499152 130898 499194 131134
rect 498874 130866 499194 130898
rect 504805 131454 505125 131486
rect 504805 131218 504847 131454
rect 505083 131218 505125 131454
rect 504805 131134 505125 131218
rect 504805 130898 504847 131134
rect 505083 130898 505125 131134
rect 504805 130866 505125 130898
rect 526874 131454 527194 131486
rect 526874 131218 526916 131454
rect 527152 131218 527194 131454
rect 526874 131134 527194 131218
rect 526874 130898 526916 131134
rect 527152 130898 527194 131134
rect 526874 130866 527194 130898
rect 532805 131454 533125 131486
rect 532805 131218 532847 131454
rect 533083 131218 533125 131454
rect 532805 131134 533125 131218
rect 532805 130898 532847 131134
rect 533083 130898 533125 131134
rect 532805 130866 533125 130898
rect 554874 131454 555194 131486
rect 554874 131218 554916 131454
rect 555152 131218 555194 131454
rect 554874 131134 555194 131218
rect 554874 130898 554916 131134
rect 555152 130898 555194 131134
rect 554874 130866 555194 130898
rect 560805 131454 561125 131486
rect 560805 131218 560847 131454
rect 561083 131218 561125 131454
rect 560805 131134 561125 131218
rect 560805 130898 560847 131134
rect 561083 130898 561125 131134
rect 560805 130866 561125 130898
rect -2006 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 -1386 107829
rect -2006 107509 -1386 107593
rect -2006 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 -1386 107509
rect -2006 80829 -1386 107273
rect 19910 107829 20230 107861
rect 19910 107593 19952 107829
rect 20188 107593 20230 107829
rect 19910 107509 20230 107593
rect 19910 107273 19952 107509
rect 20188 107273 20230 107509
rect 19910 107241 20230 107273
rect 25840 107829 26160 107861
rect 25840 107593 25882 107829
rect 26118 107593 26160 107829
rect 25840 107509 26160 107593
rect 25840 107273 25882 107509
rect 26118 107273 26160 107509
rect 25840 107241 26160 107273
rect 31771 107829 32091 107861
rect 31771 107593 31813 107829
rect 32049 107593 32091 107829
rect 31771 107509 32091 107593
rect 31771 107273 31813 107509
rect 32049 107273 32091 107509
rect 31771 107241 32091 107273
rect 47910 107829 48230 107861
rect 47910 107593 47952 107829
rect 48188 107593 48230 107829
rect 47910 107509 48230 107593
rect 47910 107273 47952 107509
rect 48188 107273 48230 107509
rect 47910 107241 48230 107273
rect 53840 107829 54160 107861
rect 53840 107593 53882 107829
rect 54118 107593 54160 107829
rect 53840 107509 54160 107593
rect 53840 107273 53882 107509
rect 54118 107273 54160 107509
rect 53840 107241 54160 107273
rect 59771 107829 60091 107861
rect 59771 107593 59813 107829
rect 60049 107593 60091 107829
rect 59771 107509 60091 107593
rect 59771 107273 59813 107509
rect 60049 107273 60091 107509
rect 59771 107241 60091 107273
rect 75910 107829 76230 107861
rect 75910 107593 75952 107829
rect 76188 107593 76230 107829
rect 75910 107509 76230 107593
rect 75910 107273 75952 107509
rect 76188 107273 76230 107509
rect 75910 107241 76230 107273
rect 81840 107829 82160 107861
rect 81840 107593 81882 107829
rect 82118 107593 82160 107829
rect 81840 107509 82160 107593
rect 81840 107273 81882 107509
rect 82118 107273 82160 107509
rect 81840 107241 82160 107273
rect 87771 107829 88091 107861
rect 87771 107593 87813 107829
rect 88049 107593 88091 107829
rect 87771 107509 88091 107593
rect 87771 107273 87813 107509
rect 88049 107273 88091 107509
rect 87771 107241 88091 107273
rect 103910 107829 104230 107861
rect 103910 107593 103952 107829
rect 104188 107593 104230 107829
rect 103910 107509 104230 107593
rect 103910 107273 103952 107509
rect 104188 107273 104230 107509
rect 103910 107241 104230 107273
rect 109840 107829 110160 107861
rect 109840 107593 109882 107829
rect 110118 107593 110160 107829
rect 109840 107509 110160 107593
rect 109840 107273 109882 107509
rect 110118 107273 110160 107509
rect 109840 107241 110160 107273
rect 115771 107829 116091 107861
rect 115771 107593 115813 107829
rect 116049 107593 116091 107829
rect 115771 107509 116091 107593
rect 115771 107273 115813 107509
rect 116049 107273 116091 107509
rect 115771 107241 116091 107273
rect 131910 107829 132230 107861
rect 131910 107593 131952 107829
rect 132188 107593 132230 107829
rect 131910 107509 132230 107593
rect 131910 107273 131952 107509
rect 132188 107273 132230 107509
rect 131910 107241 132230 107273
rect 137840 107829 138160 107861
rect 137840 107593 137882 107829
rect 138118 107593 138160 107829
rect 137840 107509 138160 107593
rect 137840 107273 137882 107509
rect 138118 107273 138160 107509
rect 137840 107241 138160 107273
rect 143771 107829 144091 107861
rect 143771 107593 143813 107829
rect 144049 107593 144091 107829
rect 143771 107509 144091 107593
rect 143771 107273 143813 107509
rect 144049 107273 144091 107509
rect 143771 107241 144091 107273
rect 159910 107829 160230 107861
rect 159910 107593 159952 107829
rect 160188 107593 160230 107829
rect 159910 107509 160230 107593
rect 159910 107273 159952 107509
rect 160188 107273 160230 107509
rect 159910 107241 160230 107273
rect 165840 107829 166160 107861
rect 165840 107593 165882 107829
rect 166118 107593 166160 107829
rect 165840 107509 166160 107593
rect 165840 107273 165882 107509
rect 166118 107273 166160 107509
rect 165840 107241 166160 107273
rect 171771 107829 172091 107861
rect 171771 107593 171813 107829
rect 172049 107593 172091 107829
rect 171771 107509 172091 107593
rect 171771 107273 171813 107509
rect 172049 107273 172091 107509
rect 171771 107241 172091 107273
rect 187910 107829 188230 107861
rect 187910 107593 187952 107829
rect 188188 107593 188230 107829
rect 187910 107509 188230 107593
rect 187910 107273 187952 107509
rect 188188 107273 188230 107509
rect 187910 107241 188230 107273
rect 193840 107829 194160 107861
rect 193840 107593 193882 107829
rect 194118 107593 194160 107829
rect 193840 107509 194160 107593
rect 193840 107273 193882 107509
rect 194118 107273 194160 107509
rect 193840 107241 194160 107273
rect 199771 107829 200091 107861
rect 199771 107593 199813 107829
rect 200049 107593 200091 107829
rect 199771 107509 200091 107593
rect 199771 107273 199813 107509
rect 200049 107273 200091 107509
rect 199771 107241 200091 107273
rect 215910 107829 216230 107861
rect 215910 107593 215952 107829
rect 216188 107593 216230 107829
rect 215910 107509 216230 107593
rect 215910 107273 215952 107509
rect 216188 107273 216230 107509
rect 215910 107241 216230 107273
rect 221840 107829 222160 107861
rect 221840 107593 221882 107829
rect 222118 107593 222160 107829
rect 221840 107509 222160 107593
rect 221840 107273 221882 107509
rect 222118 107273 222160 107509
rect 221840 107241 222160 107273
rect 227771 107829 228091 107861
rect 227771 107593 227813 107829
rect 228049 107593 228091 107829
rect 227771 107509 228091 107593
rect 227771 107273 227813 107509
rect 228049 107273 228091 107509
rect 227771 107241 228091 107273
rect 243910 107829 244230 107861
rect 243910 107593 243952 107829
rect 244188 107593 244230 107829
rect 243910 107509 244230 107593
rect 243910 107273 243952 107509
rect 244188 107273 244230 107509
rect 243910 107241 244230 107273
rect 249840 107829 250160 107861
rect 249840 107593 249882 107829
rect 250118 107593 250160 107829
rect 249840 107509 250160 107593
rect 249840 107273 249882 107509
rect 250118 107273 250160 107509
rect 249840 107241 250160 107273
rect 255771 107829 256091 107861
rect 255771 107593 255813 107829
rect 256049 107593 256091 107829
rect 255771 107509 256091 107593
rect 255771 107273 255813 107509
rect 256049 107273 256091 107509
rect 255771 107241 256091 107273
rect 271910 107829 272230 107861
rect 271910 107593 271952 107829
rect 272188 107593 272230 107829
rect 271910 107509 272230 107593
rect 271910 107273 271952 107509
rect 272188 107273 272230 107509
rect 271910 107241 272230 107273
rect 277840 107829 278160 107861
rect 277840 107593 277882 107829
rect 278118 107593 278160 107829
rect 277840 107509 278160 107593
rect 277840 107273 277882 107509
rect 278118 107273 278160 107509
rect 277840 107241 278160 107273
rect 283771 107829 284091 107861
rect 283771 107593 283813 107829
rect 284049 107593 284091 107829
rect 283771 107509 284091 107593
rect 283771 107273 283813 107509
rect 284049 107273 284091 107509
rect 283771 107241 284091 107273
rect 299910 107829 300230 107861
rect 299910 107593 299952 107829
rect 300188 107593 300230 107829
rect 299910 107509 300230 107593
rect 299910 107273 299952 107509
rect 300188 107273 300230 107509
rect 299910 107241 300230 107273
rect 305840 107829 306160 107861
rect 305840 107593 305882 107829
rect 306118 107593 306160 107829
rect 305840 107509 306160 107593
rect 305840 107273 305882 107509
rect 306118 107273 306160 107509
rect 305840 107241 306160 107273
rect 311771 107829 312091 107861
rect 311771 107593 311813 107829
rect 312049 107593 312091 107829
rect 311771 107509 312091 107593
rect 311771 107273 311813 107509
rect 312049 107273 312091 107509
rect 311771 107241 312091 107273
rect 327910 107829 328230 107861
rect 327910 107593 327952 107829
rect 328188 107593 328230 107829
rect 327910 107509 328230 107593
rect 327910 107273 327952 107509
rect 328188 107273 328230 107509
rect 327910 107241 328230 107273
rect 333840 107829 334160 107861
rect 333840 107593 333882 107829
rect 334118 107593 334160 107829
rect 333840 107509 334160 107593
rect 333840 107273 333882 107509
rect 334118 107273 334160 107509
rect 333840 107241 334160 107273
rect 339771 107829 340091 107861
rect 339771 107593 339813 107829
rect 340049 107593 340091 107829
rect 339771 107509 340091 107593
rect 339771 107273 339813 107509
rect 340049 107273 340091 107509
rect 339771 107241 340091 107273
rect 355910 107829 356230 107861
rect 355910 107593 355952 107829
rect 356188 107593 356230 107829
rect 355910 107509 356230 107593
rect 355910 107273 355952 107509
rect 356188 107273 356230 107509
rect 355910 107241 356230 107273
rect 361840 107829 362160 107861
rect 361840 107593 361882 107829
rect 362118 107593 362160 107829
rect 361840 107509 362160 107593
rect 361840 107273 361882 107509
rect 362118 107273 362160 107509
rect 361840 107241 362160 107273
rect 367771 107829 368091 107861
rect 367771 107593 367813 107829
rect 368049 107593 368091 107829
rect 367771 107509 368091 107593
rect 367771 107273 367813 107509
rect 368049 107273 368091 107509
rect 367771 107241 368091 107273
rect 383910 107829 384230 107861
rect 383910 107593 383952 107829
rect 384188 107593 384230 107829
rect 383910 107509 384230 107593
rect 383910 107273 383952 107509
rect 384188 107273 384230 107509
rect 383910 107241 384230 107273
rect 389840 107829 390160 107861
rect 389840 107593 389882 107829
rect 390118 107593 390160 107829
rect 389840 107509 390160 107593
rect 389840 107273 389882 107509
rect 390118 107273 390160 107509
rect 389840 107241 390160 107273
rect 395771 107829 396091 107861
rect 395771 107593 395813 107829
rect 396049 107593 396091 107829
rect 395771 107509 396091 107593
rect 395771 107273 395813 107509
rect 396049 107273 396091 107509
rect 395771 107241 396091 107273
rect 411910 107829 412230 107861
rect 411910 107593 411952 107829
rect 412188 107593 412230 107829
rect 411910 107509 412230 107593
rect 411910 107273 411952 107509
rect 412188 107273 412230 107509
rect 411910 107241 412230 107273
rect 417840 107829 418160 107861
rect 417840 107593 417882 107829
rect 418118 107593 418160 107829
rect 417840 107509 418160 107593
rect 417840 107273 417882 107509
rect 418118 107273 418160 107509
rect 417840 107241 418160 107273
rect 423771 107829 424091 107861
rect 423771 107593 423813 107829
rect 424049 107593 424091 107829
rect 423771 107509 424091 107593
rect 423771 107273 423813 107509
rect 424049 107273 424091 107509
rect 423771 107241 424091 107273
rect 439910 107829 440230 107861
rect 439910 107593 439952 107829
rect 440188 107593 440230 107829
rect 439910 107509 440230 107593
rect 439910 107273 439952 107509
rect 440188 107273 440230 107509
rect 439910 107241 440230 107273
rect 445840 107829 446160 107861
rect 445840 107593 445882 107829
rect 446118 107593 446160 107829
rect 445840 107509 446160 107593
rect 445840 107273 445882 107509
rect 446118 107273 446160 107509
rect 445840 107241 446160 107273
rect 451771 107829 452091 107861
rect 451771 107593 451813 107829
rect 452049 107593 452091 107829
rect 451771 107509 452091 107593
rect 451771 107273 451813 107509
rect 452049 107273 452091 107509
rect 451771 107241 452091 107273
rect 467910 107829 468230 107861
rect 467910 107593 467952 107829
rect 468188 107593 468230 107829
rect 467910 107509 468230 107593
rect 467910 107273 467952 107509
rect 468188 107273 468230 107509
rect 467910 107241 468230 107273
rect 473840 107829 474160 107861
rect 473840 107593 473882 107829
rect 474118 107593 474160 107829
rect 473840 107509 474160 107593
rect 473840 107273 473882 107509
rect 474118 107273 474160 107509
rect 473840 107241 474160 107273
rect 479771 107829 480091 107861
rect 479771 107593 479813 107829
rect 480049 107593 480091 107829
rect 479771 107509 480091 107593
rect 479771 107273 479813 107509
rect 480049 107273 480091 107509
rect 479771 107241 480091 107273
rect 495910 107829 496230 107861
rect 495910 107593 495952 107829
rect 496188 107593 496230 107829
rect 495910 107509 496230 107593
rect 495910 107273 495952 107509
rect 496188 107273 496230 107509
rect 495910 107241 496230 107273
rect 501840 107829 502160 107861
rect 501840 107593 501882 107829
rect 502118 107593 502160 107829
rect 501840 107509 502160 107593
rect 501840 107273 501882 107509
rect 502118 107273 502160 107509
rect 501840 107241 502160 107273
rect 507771 107829 508091 107861
rect 507771 107593 507813 107829
rect 508049 107593 508091 107829
rect 507771 107509 508091 107593
rect 507771 107273 507813 107509
rect 508049 107273 508091 107509
rect 507771 107241 508091 107273
rect 523910 107829 524230 107861
rect 523910 107593 523952 107829
rect 524188 107593 524230 107829
rect 523910 107509 524230 107593
rect 523910 107273 523952 107509
rect 524188 107273 524230 107509
rect 523910 107241 524230 107273
rect 529840 107829 530160 107861
rect 529840 107593 529882 107829
rect 530118 107593 530160 107829
rect 529840 107509 530160 107593
rect 529840 107273 529882 107509
rect 530118 107273 530160 107509
rect 529840 107241 530160 107273
rect 535771 107829 536091 107861
rect 535771 107593 535813 107829
rect 536049 107593 536091 107829
rect 535771 107509 536091 107593
rect 535771 107273 535813 107509
rect 536049 107273 536091 107509
rect 535771 107241 536091 107273
rect 551910 107829 552230 107861
rect 551910 107593 551952 107829
rect 552188 107593 552230 107829
rect 551910 107509 552230 107593
rect 551910 107273 551952 107509
rect 552188 107273 552230 107509
rect 551910 107241 552230 107273
rect 557840 107829 558160 107861
rect 557840 107593 557882 107829
rect 558118 107593 558160 107829
rect 557840 107509 558160 107593
rect 557840 107273 557882 107509
rect 558118 107273 558160 107509
rect 557840 107241 558160 107273
rect 563771 107829 564091 107861
rect 563771 107593 563813 107829
rect 564049 107593 564091 107829
rect 563771 107509 564091 107593
rect 563771 107273 563813 107509
rect 564049 107273 564091 107509
rect 563771 107241 564091 107273
rect 573494 107829 574114 134273
rect 573494 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 574114 107829
rect 573494 107509 574114 107593
rect 573494 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 574114 107509
rect 22874 104454 23194 104486
rect 22874 104218 22916 104454
rect 23152 104218 23194 104454
rect 22874 104134 23194 104218
rect 22874 103898 22916 104134
rect 23152 103898 23194 104134
rect 22874 103866 23194 103898
rect 28805 104454 29125 104486
rect 28805 104218 28847 104454
rect 29083 104218 29125 104454
rect 28805 104134 29125 104218
rect 28805 103898 28847 104134
rect 29083 103898 29125 104134
rect 28805 103866 29125 103898
rect 50874 104454 51194 104486
rect 50874 104218 50916 104454
rect 51152 104218 51194 104454
rect 50874 104134 51194 104218
rect 50874 103898 50916 104134
rect 51152 103898 51194 104134
rect 50874 103866 51194 103898
rect 56805 104454 57125 104486
rect 56805 104218 56847 104454
rect 57083 104218 57125 104454
rect 56805 104134 57125 104218
rect 56805 103898 56847 104134
rect 57083 103898 57125 104134
rect 56805 103866 57125 103898
rect 78874 104454 79194 104486
rect 78874 104218 78916 104454
rect 79152 104218 79194 104454
rect 78874 104134 79194 104218
rect 78874 103898 78916 104134
rect 79152 103898 79194 104134
rect 78874 103866 79194 103898
rect 84805 104454 85125 104486
rect 84805 104218 84847 104454
rect 85083 104218 85125 104454
rect 84805 104134 85125 104218
rect 84805 103898 84847 104134
rect 85083 103898 85125 104134
rect 84805 103866 85125 103898
rect 106874 104454 107194 104486
rect 106874 104218 106916 104454
rect 107152 104218 107194 104454
rect 106874 104134 107194 104218
rect 106874 103898 106916 104134
rect 107152 103898 107194 104134
rect 106874 103866 107194 103898
rect 112805 104454 113125 104486
rect 112805 104218 112847 104454
rect 113083 104218 113125 104454
rect 112805 104134 113125 104218
rect 112805 103898 112847 104134
rect 113083 103898 113125 104134
rect 112805 103866 113125 103898
rect 134874 104454 135194 104486
rect 134874 104218 134916 104454
rect 135152 104218 135194 104454
rect 134874 104134 135194 104218
rect 134874 103898 134916 104134
rect 135152 103898 135194 104134
rect 134874 103866 135194 103898
rect 140805 104454 141125 104486
rect 140805 104218 140847 104454
rect 141083 104218 141125 104454
rect 140805 104134 141125 104218
rect 140805 103898 140847 104134
rect 141083 103898 141125 104134
rect 140805 103866 141125 103898
rect 162874 104454 163194 104486
rect 162874 104218 162916 104454
rect 163152 104218 163194 104454
rect 162874 104134 163194 104218
rect 162874 103898 162916 104134
rect 163152 103898 163194 104134
rect 162874 103866 163194 103898
rect 168805 104454 169125 104486
rect 168805 104218 168847 104454
rect 169083 104218 169125 104454
rect 168805 104134 169125 104218
rect 168805 103898 168847 104134
rect 169083 103898 169125 104134
rect 168805 103866 169125 103898
rect 190874 104454 191194 104486
rect 190874 104218 190916 104454
rect 191152 104218 191194 104454
rect 190874 104134 191194 104218
rect 190874 103898 190916 104134
rect 191152 103898 191194 104134
rect 190874 103866 191194 103898
rect 196805 104454 197125 104486
rect 196805 104218 196847 104454
rect 197083 104218 197125 104454
rect 196805 104134 197125 104218
rect 196805 103898 196847 104134
rect 197083 103898 197125 104134
rect 196805 103866 197125 103898
rect 218874 104454 219194 104486
rect 218874 104218 218916 104454
rect 219152 104218 219194 104454
rect 218874 104134 219194 104218
rect 218874 103898 218916 104134
rect 219152 103898 219194 104134
rect 218874 103866 219194 103898
rect 224805 104454 225125 104486
rect 224805 104218 224847 104454
rect 225083 104218 225125 104454
rect 224805 104134 225125 104218
rect 224805 103898 224847 104134
rect 225083 103898 225125 104134
rect 224805 103866 225125 103898
rect 246874 104454 247194 104486
rect 246874 104218 246916 104454
rect 247152 104218 247194 104454
rect 246874 104134 247194 104218
rect 246874 103898 246916 104134
rect 247152 103898 247194 104134
rect 246874 103866 247194 103898
rect 252805 104454 253125 104486
rect 252805 104218 252847 104454
rect 253083 104218 253125 104454
rect 252805 104134 253125 104218
rect 252805 103898 252847 104134
rect 253083 103898 253125 104134
rect 252805 103866 253125 103898
rect 274874 104454 275194 104486
rect 274874 104218 274916 104454
rect 275152 104218 275194 104454
rect 274874 104134 275194 104218
rect 274874 103898 274916 104134
rect 275152 103898 275194 104134
rect 274874 103866 275194 103898
rect 280805 104454 281125 104486
rect 280805 104218 280847 104454
rect 281083 104218 281125 104454
rect 280805 104134 281125 104218
rect 280805 103898 280847 104134
rect 281083 103898 281125 104134
rect 280805 103866 281125 103898
rect 302874 104454 303194 104486
rect 302874 104218 302916 104454
rect 303152 104218 303194 104454
rect 302874 104134 303194 104218
rect 302874 103898 302916 104134
rect 303152 103898 303194 104134
rect 302874 103866 303194 103898
rect 308805 104454 309125 104486
rect 308805 104218 308847 104454
rect 309083 104218 309125 104454
rect 308805 104134 309125 104218
rect 308805 103898 308847 104134
rect 309083 103898 309125 104134
rect 308805 103866 309125 103898
rect 330874 104454 331194 104486
rect 330874 104218 330916 104454
rect 331152 104218 331194 104454
rect 330874 104134 331194 104218
rect 330874 103898 330916 104134
rect 331152 103898 331194 104134
rect 330874 103866 331194 103898
rect 336805 104454 337125 104486
rect 336805 104218 336847 104454
rect 337083 104218 337125 104454
rect 336805 104134 337125 104218
rect 336805 103898 336847 104134
rect 337083 103898 337125 104134
rect 336805 103866 337125 103898
rect 358874 104454 359194 104486
rect 358874 104218 358916 104454
rect 359152 104218 359194 104454
rect 358874 104134 359194 104218
rect 358874 103898 358916 104134
rect 359152 103898 359194 104134
rect 358874 103866 359194 103898
rect 364805 104454 365125 104486
rect 364805 104218 364847 104454
rect 365083 104218 365125 104454
rect 364805 104134 365125 104218
rect 364805 103898 364847 104134
rect 365083 103898 365125 104134
rect 364805 103866 365125 103898
rect 386874 104454 387194 104486
rect 386874 104218 386916 104454
rect 387152 104218 387194 104454
rect 386874 104134 387194 104218
rect 386874 103898 386916 104134
rect 387152 103898 387194 104134
rect 386874 103866 387194 103898
rect 392805 104454 393125 104486
rect 392805 104218 392847 104454
rect 393083 104218 393125 104454
rect 392805 104134 393125 104218
rect 392805 103898 392847 104134
rect 393083 103898 393125 104134
rect 392805 103866 393125 103898
rect 414874 104454 415194 104486
rect 414874 104218 414916 104454
rect 415152 104218 415194 104454
rect 414874 104134 415194 104218
rect 414874 103898 414916 104134
rect 415152 103898 415194 104134
rect 414874 103866 415194 103898
rect 420805 104454 421125 104486
rect 420805 104218 420847 104454
rect 421083 104218 421125 104454
rect 420805 104134 421125 104218
rect 420805 103898 420847 104134
rect 421083 103898 421125 104134
rect 420805 103866 421125 103898
rect 442874 104454 443194 104486
rect 442874 104218 442916 104454
rect 443152 104218 443194 104454
rect 442874 104134 443194 104218
rect 442874 103898 442916 104134
rect 443152 103898 443194 104134
rect 442874 103866 443194 103898
rect 448805 104454 449125 104486
rect 448805 104218 448847 104454
rect 449083 104218 449125 104454
rect 448805 104134 449125 104218
rect 448805 103898 448847 104134
rect 449083 103898 449125 104134
rect 448805 103866 449125 103898
rect 470874 104454 471194 104486
rect 470874 104218 470916 104454
rect 471152 104218 471194 104454
rect 470874 104134 471194 104218
rect 470874 103898 470916 104134
rect 471152 103898 471194 104134
rect 470874 103866 471194 103898
rect 476805 104454 477125 104486
rect 476805 104218 476847 104454
rect 477083 104218 477125 104454
rect 476805 104134 477125 104218
rect 476805 103898 476847 104134
rect 477083 103898 477125 104134
rect 476805 103866 477125 103898
rect 498874 104454 499194 104486
rect 498874 104218 498916 104454
rect 499152 104218 499194 104454
rect 498874 104134 499194 104218
rect 498874 103898 498916 104134
rect 499152 103898 499194 104134
rect 498874 103866 499194 103898
rect 504805 104454 505125 104486
rect 504805 104218 504847 104454
rect 505083 104218 505125 104454
rect 504805 104134 505125 104218
rect 504805 103898 504847 104134
rect 505083 103898 505125 104134
rect 504805 103866 505125 103898
rect 526874 104454 527194 104486
rect 526874 104218 526916 104454
rect 527152 104218 527194 104454
rect 526874 104134 527194 104218
rect 526874 103898 526916 104134
rect 527152 103898 527194 104134
rect 526874 103866 527194 103898
rect 532805 104454 533125 104486
rect 532805 104218 532847 104454
rect 533083 104218 533125 104454
rect 532805 104134 533125 104218
rect 532805 103898 532847 104134
rect 533083 103898 533125 104134
rect 532805 103866 533125 103898
rect 554874 104454 555194 104486
rect 554874 104218 554916 104454
rect 555152 104218 555194 104454
rect 554874 104134 555194 104218
rect 554874 103898 554916 104134
rect 555152 103898 555194 104134
rect 554874 103866 555194 103898
rect 560805 104454 561125 104486
rect 560805 104218 560847 104454
rect 561083 104218 561125 104454
rect 560805 104134 561125 104218
rect 560805 103898 560847 104134
rect 561083 103898 561125 104134
rect 560805 103866 561125 103898
rect -2006 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 -1386 80829
rect -2006 80509 -1386 80593
rect -2006 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 -1386 80509
rect -2006 53829 -1386 80273
rect 19910 80829 20230 80861
rect 19910 80593 19952 80829
rect 20188 80593 20230 80829
rect 19910 80509 20230 80593
rect 19910 80273 19952 80509
rect 20188 80273 20230 80509
rect 19910 80241 20230 80273
rect 25840 80829 26160 80861
rect 25840 80593 25882 80829
rect 26118 80593 26160 80829
rect 25840 80509 26160 80593
rect 25840 80273 25882 80509
rect 26118 80273 26160 80509
rect 25840 80241 26160 80273
rect 31771 80829 32091 80861
rect 31771 80593 31813 80829
rect 32049 80593 32091 80829
rect 31771 80509 32091 80593
rect 31771 80273 31813 80509
rect 32049 80273 32091 80509
rect 31771 80241 32091 80273
rect 47910 80829 48230 80861
rect 47910 80593 47952 80829
rect 48188 80593 48230 80829
rect 47910 80509 48230 80593
rect 47910 80273 47952 80509
rect 48188 80273 48230 80509
rect 47910 80241 48230 80273
rect 53840 80829 54160 80861
rect 53840 80593 53882 80829
rect 54118 80593 54160 80829
rect 53840 80509 54160 80593
rect 53840 80273 53882 80509
rect 54118 80273 54160 80509
rect 53840 80241 54160 80273
rect 59771 80829 60091 80861
rect 59771 80593 59813 80829
rect 60049 80593 60091 80829
rect 59771 80509 60091 80593
rect 59771 80273 59813 80509
rect 60049 80273 60091 80509
rect 59771 80241 60091 80273
rect 75910 80829 76230 80861
rect 75910 80593 75952 80829
rect 76188 80593 76230 80829
rect 75910 80509 76230 80593
rect 75910 80273 75952 80509
rect 76188 80273 76230 80509
rect 75910 80241 76230 80273
rect 81840 80829 82160 80861
rect 81840 80593 81882 80829
rect 82118 80593 82160 80829
rect 81840 80509 82160 80593
rect 81840 80273 81882 80509
rect 82118 80273 82160 80509
rect 81840 80241 82160 80273
rect 87771 80829 88091 80861
rect 87771 80593 87813 80829
rect 88049 80593 88091 80829
rect 87771 80509 88091 80593
rect 87771 80273 87813 80509
rect 88049 80273 88091 80509
rect 87771 80241 88091 80273
rect 103910 80829 104230 80861
rect 103910 80593 103952 80829
rect 104188 80593 104230 80829
rect 103910 80509 104230 80593
rect 103910 80273 103952 80509
rect 104188 80273 104230 80509
rect 103910 80241 104230 80273
rect 109840 80829 110160 80861
rect 109840 80593 109882 80829
rect 110118 80593 110160 80829
rect 109840 80509 110160 80593
rect 109840 80273 109882 80509
rect 110118 80273 110160 80509
rect 109840 80241 110160 80273
rect 115771 80829 116091 80861
rect 115771 80593 115813 80829
rect 116049 80593 116091 80829
rect 115771 80509 116091 80593
rect 115771 80273 115813 80509
rect 116049 80273 116091 80509
rect 115771 80241 116091 80273
rect 131910 80829 132230 80861
rect 131910 80593 131952 80829
rect 132188 80593 132230 80829
rect 131910 80509 132230 80593
rect 131910 80273 131952 80509
rect 132188 80273 132230 80509
rect 131910 80241 132230 80273
rect 137840 80829 138160 80861
rect 137840 80593 137882 80829
rect 138118 80593 138160 80829
rect 137840 80509 138160 80593
rect 137840 80273 137882 80509
rect 138118 80273 138160 80509
rect 137840 80241 138160 80273
rect 143771 80829 144091 80861
rect 143771 80593 143813 80829
rect 144049 80593 144091 80829
rect 143771 80509 144091 80593
rect 143771 80273 143813 80509
rect 144049 80273 144091 80509
rect 143771 80241 144091 80273
rect 159910 80829 160230 80861
rect 159910 80593 159952 80829
rect 160188 80593 160230 80829
rect 159910 80509 160230 80593
rect 159910 80273 159952 80509
rect 160188 80273 160230 80509
rect 159910 80241 160230 80273
rect 165840 80829 166160 80861
rect 165840 80593 165882 80829
rect 166118 80593 166160 80829
rect 165840 80509 166160 80593
rect 165840 80273 165882 80509
rect 166118 80273 166160 80509
rect 165840 80241 166160 80273
rect 171771 80829 172091 80861
rect 171771 80593 171813 80829
rect 172049 80593 172091 80829
rect 171771 80509 172091 80593
rect 171771 80273 171813 80509
rect 172049 80273 172091 80509
rect 171771 80241 172091 80273
rect 187910 80829 188230 80861
rect 187910 80593 187952 80829
rect 188188 80593 188230 80829
rect 187910 80509 188230 80593
rect 187910 80273 187952 80509
rect 188188 80273 188230 80509
rect 187910 80241 188230 80273
rect 193840 80829 194160 80861
rect 193840 80593 193882 80829
rect 194118 80593 194160 80829
rect 193840 80509 194160 80593
rect 193840 80273 193882 80509
rect 194118 80273 194160 80509
rect 193840 80241 194160 80273
rect 199771 80829 200091 80861
rect 199771 80593 199813 80829
rect 200049 80593 200091 80829
rect 199771 80509 200091 80593
rect 199771 80273 199813 80509
rect 200049 80273 200091 80509
rect 199771 80241 200091 80273
rect 215910 80829 216230 80861
rect 215910 80593 215952 80829
rect 216188 80593 216230 80829
rect 215910 80509 216230 80593
rect 215910 80273 215952 80509
rect 216188 80273 216230 80509
rect 215910 80241 216230 80273
rect 221840 80829 222160 80861
rect 221840 80593 221882 80829
rect 222118 80593 222160 80829
rect 221840 80509 222160 80593
rect 221840 80273 221882 80509
rect 222118 80273 222160 80509
rect 221840 80241 222160 80273
rect 227771 80829 228091 80861
rect 227771 80593 227813 80829
rect 228049 80593 228091 80829
rect 227771 80509 228091 80593
rect 227771 80273 227813 80509
rect 228049 80273 228091 80509
rect 227771 80241 228091 80273
rect 243910 80829 244230 80861
rect 243910 80593 243952 80829
rect 244188 80593 244230 80829
rect 243910 80509 244230 80593
rect 243910 80273 243952 80509
rect 244188 80273 244230 80509
rect 243910 80241 244230 80273
rect 249840 80829 250160 80861
rect 249840 80593 249882 80829
rect 250118 80593 250160 80829
rect 249840 80509 250160 80593
rect 249840 80273 249882 80509
rect 250118 80273 250160 80509
rect 249840 80241 250160 80273
rect 255771 80829 256091 80861
rect 255771 80593 255813 80829
rect 256049 80593 256091 80829
rect 255771 80509 256091 80593
rect 255771 80273 255813 80509
rect 256049 80273 256091 80509
rect 255771 80241 256091 80273
rect 271910 80829 272230 80861
rect 271910 80593 271952 80829
rect 272188 80593 272230 80829
rect 271910 80509 272230 80593
rect 271910 80273 271952 80509
rect 272188 80273 272230 80509
rect 271910 80241 272230 80273
rect 277840 80829 278160 80861
rect 277840 80593 277882 80829
rect 278118 80593 278160 80829
rect 277840 80509 278160 80593
rect 277840 80273 277882 80509
rect 278118 80273 278160 80509
rect 277840 80241 278160 80273
rect 283771 80829 284091 80861
rect 283771 80593 283813 80829
rect 284049 80593 284091 80829
rect 283771 80509 284091 80593
rect 283771 80273 283813 80509
rect 284049 80273 284091 80509
rect 283771 80241 284091 80273
rect 299910 80829 300230 80861
rect 299910 80593 299952 80829
rect 300188 80593 300230 80829
rect 299910 80509 300230 80593
rect 299910 80273 299952 80509
rect 300188 80273 300230 80509
rect 299910 80241 300230 80273
rect 305840 80829 306160 80861
rect 305840 80593 305882 80829
rect 306118 80593 306160 80829
rect 305840 80509 306160 80593
rect 305840 80273 305882 80509
rect 306118 80273 306160 80509
rect 305840 80241 306160 80273
rect 311771 80829 312091 80861
rect 311771 80593 311813 80829
rect 312049 80593 312091 80829
rect 311771 80509 312091 80593
rect 311771 80273 311813 80509
rect 312049 80273 312091 80509
rect 311771 80241 312091 80273
rect 327910 80829 328230 80861
rect 327910 80593 327952 80829
rect 328188 80593 328230 80829
rect 327910 80509 328230 80593
rect 327910 80273 327952 80509
rect 328188 80273 328230 80509
rect 327910 80241 328230 80273
rect 333840 80829 334160 80861
rect 333840 80593 333882 80829
rect 334118 80593 334160 80829
rect 333840 80509 334160 80593
rect 333840 80273 333882 80509
rect 334118 80273 334160 80509
rect 333840 80241 334160 80273
rect 339771 80829 340091 80861
rect 339771 80593 339813 80829
rect 340049 80593 340091 80829
rect 339771 80509 340091 80593
rect 339771 80273 339813 80509
rect 340049 80273 340091 80509
rect 339771 80241 340091 80273
rect 355910 80829 356230 80861
rect 355910 80593 355952 80829
rect 356188 80593 356230 80829
rect 355910 80509 356230 80593
rect 355910 80273 355952 80509
rect 356188 80273 356230 80509
rect 355910 80241 356230 80273
rect 361840 80829 362160 80861
rect 361840 80593 361882 80829
rect 362118 80593 362160 80829
rect 361840 80509 362160 80593
rect 361840 80273 361882 80509
rect 362118 80273 362160 80509
rect 361840 80241 362160 80273
rect 367771 80829 368091 80861
rect 367771 80593 367813 80829
rect 368049 80593 368091 80829
rect 367771 80509 368091 80593
rect 367771 80273 367813 80509
rect 368049 80273 368091 80509
rect 367771 80241 368091 80273
rect 383910 80829 384230 80861
rect 383910 80593 383952 80829
rect 384188 80593 384230 80829
rect 383910 80509 384230 80593
rect 383910 80273 383952 80509
rect 384188 80273 384230 80509
rect 383910 80241 384230 80273
rect 389840 80829 390160 80861
rect 389840 80593 389882 80829
rect 390118 80593 390160 80829
rect 389840 80509 390160 80593
rect 389840 80273 389882 80509
rect 390118 80273 390160 80509
rect 389840 80241 390160 80273
rect 395771 80829 396091 80861
rect 395771 80593 395813 80829
rect 396049 80593 396091 80829
rect 395771 80509 396091 80593
rect 395771 80273 395813 80509
rect 396049 80273 396091 80509
rect 395771 80241 396091 80273
rect 411910 80829 412230 80861
rect 411910 80593 411952 80829
rect 412188 80593 412230 80829
rect 411910 80509 412230 80593
rect 411910 80273 411952 80509
rect 412188 80273 412230 80509
rect 411910 80241 412230 80273
rect 417840 80829 418160 80861
rect 417840 80593 417882 80829
rect 418118 80593 418160 80829
rect 417840 80509 418160 80593
rect 417840 80273 417882 80509
rect 418118 80273 418160 80509
rect 417840 80241 418160 80273
rect 423771 80829 424091 80861
rect 423771 80593 423813 80829
rect 424049 80593 424091 80829
rect 423771 80509 424091 80593
rect 423771 80273 423813 80509
rect 424049 80273 424091 80509
rect 423771 80241 424091 80273
rect 439910 80829 440230 80861
rect 439910 80593 439952 80829
rect 440188 80593 440230 80829
rect 439910 80509 440230 80593
rect 439910 80273 439952 80509
rect 440188 80273 440230 80509
rect 439910 80241 440230 80273
rect 445840 80829 446160 80861
rect 445840 80593 445882 80829
rect 446118 80593 446160 80829
rect 445840 80509 446160 80593
rect 445840 80273 445882 80509
rect 446118 80273 446160 80509
rect 445840 80241 446160 80273
rect 451771 80829 452091 80861
rect 451771 80593 451813 80829
rect 452049 80593 452091 80829
rect 451771 80509 452091 80593
rect 451771 80273 451813 80509
rect 452049 80273 452091 80509
rect 451771 80241 452091 80273
rect 467910 80829 468230 80861
rect 467910 80593 467952 80829
rect 468188 80593 468230 80829
rect 467910 80509 468230 80593
rect 467910 80273 467952 80509
rect 468188 80273 468230 80509
rect 467910 80241 468230 80273
rect 473840 80829 474160 80861
rect 473840 80593 473882 80829
rect 474118 80593 474160 80829
rect 473840 80509 474160 80593
rect 473840 80273 473882 80509
rect 474118 80273 474160 80509
rect 473840 80241 474160 80273
rect 479771 80829 480091 80861
rect 479771 80593 479813 80829
rect 480049 80593 480091 80829
rect 479771 80509 480091 80593
rect 479771 80273 479813 80509
rect 480049 80273 480091 80509
rect 479771 80241 480091 80273
rect 495910 80829 496230 80861
rect 495910 80593 495952 80829
rect 496188 80593 496230 80829
rect 495910 80509 496230 80593
rect 495910 80273 495952 80509
rect 496188 80273 496230 80509
rect 495910 80241 496230 80273
rect 501840 80829 502160 80861
rect 501840 80593 501882 80829
rect 502118 80593 502160 80829
rect 501840 80509 502160 80593
rect 501840 80273 501882 80509
rect 502118 80273 502160 80509
rect 501840 80241 502160 80273
rect 507771 80829 508091 80861
rect 507771 80593 507813 80829
rect 508049 80593 508091 80829
rect 507771 80509 508091 80593
rect 507771 80273 507813 80509
rect 508049 80273 508091 80509
rect 507771 80241 508091 80273
rect 523910 80829 524230 80861
rect 523910 80593 523952 80829
rect 524188 80593 524230 80829
rect 523910 80509 524230 80593
rect 523910 80273 523952 80509
rect 524188 80273 524230 80509
rect 523910 80241 524230 80273
rect 529840 80829 530160 80861
rect 529840 80593 529882 80829
rect 530118 80593 530160 80829
rect 529840 80509 530160 80593
rect 529840 80273 529882 80509
rect 530118 80273 530160 80509
rect 529840 80241 530160 80273
rect 535771 80829 536091 80861
rect 535771 80593 535813 80829
rect 536049 80593 536091 80829
rect 535771 80509 536091 80593
rect 535771 80273 535813 80509
rect 536049 80273 536091 80509
rect 535771 80241 536091 80273
rect 551910 80829 552230 80861
rect 551910 80593 551952 80829
rect 552188 80593 552230 80829
rect 551910 80509 552230 80593
rect 551910 80273 551952 80509
rect 552188 80273 552230 80509
rect 551910 80241 552230 80273
rect 557840 80829 558160 80861
rect 557840 80593 557882 80829
rect 558118 80593 558160 80829
rect 557840 80509 558160 80593
rect 557840 80273 557882 80509
rect 558118 80273 558160 80509
rect 557840 80241 558160 80273
rect 563771 80829 564091 80861
rect 563771 80593 563813 80829
rect 564049 80593 564091 80829
rect 563771 80509 564091 80593
rect 563771 80273 563813 80509
rect 564049 80273 564091 80509
rect 563771 80241 564091 80273
rect 573494 80829 574114 107273
rect 573494 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 574114 80829
rect 573494 80509 574114 80593
rect 573494 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 574114 80509
rect 22874 77454 23194 77486
rect 22874 77218 22916 77454
rect 23152 77218 23194 77454
rect 22874 77134 23194 77218
rect 22874 76898 22916 77134
rect 23152 76898 23194 77134
rect 22874 76866 23194 76898
rect 28805 77454 29125 77486
rect 28805 77218 28847 77454
rect 29083 77218 29125 77454
rect 28805 77134 29125 77218
rect 28805 76898 28847 77134
rect 29083 76898 29125 77134
rect 28805 76866 29125 76898
rect 50874 77454 51194 77486
rect 50874 77218 50916 77454
rect 51152 77218 51194 77454
rect 50874 77134 51194 77218
rect 50874 76898 50916 77134
rect 51152 76898 51194 77134
rect 50874 76866 51194 76898
rect 56805 77454 57125 77486
rect 56805 77218 56847 77454
rect 57083 77218 57125 77454
rect 56805 77134 57125 77218
rect 56805 76898 56847 77134
rect 57083 76898 57125 77134
rect 56805 76866 57125 76898
rect 78874 77454 79194 77486
rect 78874 77218 78916 77454
rect 79152 77218 79194 77454
rect 78874 77134 79194 77218
rect 78874 76898 78916 77134
rect 79152 76898 79194 77134
rect 78874 76866 79194 76898
rect 84805 77454 85125 77486
rect 84805 77218 84847 77454
rect 85083 77218 85125 77454
rect 84805 77134 85125 77218
rect 84805 76898 84847 77134
rect 85083 76898 85125 77134
rect 84805 76866 85125 76898
rect 106874 77454 107194 77486
rect 106874 77218 106916 77454
rect 107152 77218 107194 77454
rect 106874 77134 107194 77218
rect 106874 76898 106916 77134
rect 107152 76898 107194 77134
rect 106874 76866 107194 76898
rect 112805 77454 113125 77486
rect 112805 77218 112847 77454
rect 113083 77218 113125 77454
rect 112805 77134 113125 77218
rect 112805 76898 112847 77134
rect 113083 76898 113125 77134
rect 112805 76866 113125 76898
rect 134874 77454 135194 77486
rect 134874 77218 134916 77454
rect 135152 77218 135194 77454
rect 134874 77134 135194 77218
rect 134874 76898 134916 77134
rect 135152 76898 135194 77134
rect 134874 76866 135194 76898
rect 140805 77454 141125 77486
rect 140805 77218 140847 77454
rect 141083 77218 141125 77454
rect 140805 77134 141125 77218
rect 140805 76898 140847 77134
rect 141083 76898 141125 77134
rect 140805 76866 141125 76898
rect 162874 77454 163194 77486
rect 162874 77218 162916 77454
rect 163152 77218 163194 77454
rect 162874 77134 163194 77218
rect 162874 76898 162916 77134
rect 163152 76898 163194 77134
rect 162874 76866 163194 76898
rect 168805 77454 169125 77486
rect 168805 77218 168847 77454
rect 169083 77218 169125 77454
rect 168805 77134 169125 77218
rect 168805 76898 168847 77134
rect 169083 76898 169125 77134
rect 168805 76866 169125 76898
rect 190874 77454 191194 77486
rect 190874 77218 190916 77454
rect 191152 77218 191194 77454
rect 190874 77134 191194 77218
rect 190874 76898 190916 77134
rect 191152 76898 191194 77134
rect 190874 76866 191194 76898
rect 196805 77454 197125 77486
rect 196805 77218 196847 77454
rect 197083 77218 197125 77454
rect 196805 77134 197125 77218
rect 196805 76898 196847 77134
rect 197083 76898 197125 77134
rect 196805 76866 197125 76898
rect 218874 77454 219194 77486
rect 218874 77218 218916 77454
rect 219152 77218 219194 77454
rect 218874 77134 219194 77218
rect 218874 76898 218916 77134
rect 219152 76898 219194 77134
rect 218874 76866 219194 76898
rect 224805 77454 225125 77486
rect 224805 77218 224847 77454
rect 225083 77218 225125 77454
rect 224805 77134 225125 77218
rect 224805 76898 224847 77134
rect 225083 76898 225125 77134
rect 224805 76866 225125 76898
rect 246874 77454 247194 77486
rect 246874 77218 246916 77454
rect 247152 77218 247194 77454
rect 246874 77134 247194 77218
rect 246874 76898 246916 77134
rect 247152 76898 247194 77134
rect 246874 76866 247194 76898
rect 252805 77454 253125 77486
rect 252805 77218 252847 77454
rect 253083 77218 253125 77454
rect 252805 77134 253125 77218
rect 252805 76898 252847 77134
rect 253083 76898 253125 77134
rect 252805 76866 253125 76898
rect 274874 77454 275194 77486
rect 274874 77218 274916 77454
rect 275152 77218 275194 77454
rect 274874 77134 275194 77218
rect 274874 76898 274916 77134
rect 275152 76898 275194 77134
rect 274874 76866 275194 76898
rect 280805 77454 281125 77486
rect 280805 77218 280847 77454
rect 281083 77218 281125 77454
rect 280805 77134 281125 77218
rect 280805 76898 280847 77134
rect 281083 76898 281125 77134
rect 280805 76866 281125 76898
rect 302874 77454 303194 77486
rect 302874 77218 302916 77454
rect 303152 77218 303194 77454
rect 302874 77134 303194 77218
rect 302874 76898 302916 77134
rect 303152 76898 303194 77134
rect 302874 76866 303194 76898
rect 308805 77454 309125 77486
rect 308805 77218 308847 77454
rect 309083 77218 309125 77454
rect 308805 77134 309125 77218
rect 308805 76898 308847 77134
rect 309083 76898 309125 77134
rect 308805 76866 309125 76898
rect 330874 77454 331194 77486
rect 330874 77218 330916 77454
rect 331152 77218 331194 77454
rect 330874 77134 331194 77218
rect 330874 76898 330916 77134
rect 331152 76898 331194 77134
rect 330874 76866 331194 76898
rect 336805 77454 337125 77486
rect 336805 77218 336847 77454
rect 337083 77218 337125 77454
rect 336805 77134 337125 77218
rect 336805 76898 336847 77134
rect 337083 76898 337125 77134
rect 336805 76866 337125 76898
rect 358874 77454 359194 77486
rect 358874 77218 358916 77454
rect 359152 77218 359194 77454
rect 358874 77134 359194 77218
rect 358874 76898 358916 77134
rect 359152 76898 359194 77134
rect 358874 76866 359194 76898
rect 364805 77454 365125 77486
rect 364805 77218 364847 77454
rect 365083 77218 365125 77454
rect 364805 77134 365125 77218
rect 364805 76898 364847 77134
rect 365083 76898 365125 77134
rect 364805 76866 365125 76898
rect 386874 77454 387194 77486
rect 386874 77218 386916 77454
rect 387152 77218 387194 77454
rect 386874 77134 387194 77218
rect 386874 76898 386916 77134
rect 387152 76898 387194 77134
rect 386874 76866 387194 76898
rect 392805 77454 393125 77486
rect 392805 77218 392847 77454
rect 393083 77218 393125 77454
rect 392805 77134 393125 77218
rect 392805 76898 392847 77134
rect 393083 76898 393125 77134
rect 392805 76866 393125 76898
rect 414874 77454 415194 77486
rect 414874 77218 414916 77454
rect 415152 77218 415194 77454
rect 414874 77134 415194 77218
rect 414874 76898 414916 77134
rect 415152 76898 415194 77134
rect 414874 76866 415194 76898
rect 420805 77454 421125 77486
rect 420805 77218 420847 77454
rect 421083 77218 421125 77454
rect 420805 77134 421125 77218
rect 420805 76898 420847 77134
rect 421083 76898 421125 77134
rect 420805 76866 421125 76898
rect 442874 77454 443194 77486
rect 442874 77218 442916 77454
rect 443152 77218 443194 77454
rect 442874 77134 443194 77218
rect 442874 76898 442916 77134
rect 443152 76898 443194 77134
rect 442874 76866 443194 76898
rect 448805 77454 449125 77486
rect 448805 77218 448847 77454
rect 449083 77218 449125 77454
rect 448805 77134 449125 77218
rect 448805 76898 448847 77134
rect 449083 76898 449125 77134
rect 448805 76866 449125 76898
rect 470874 77454 471194 77486
rect 470874 77218 470916 77454
rect 471152 77218 471194 77454
rect 470874 77134 471194 77218
rect 470874 76898 470916 77134
rect 471152 76898 471194 77134
rect 470874 76866 471194 76898
rect 476805 77454 477125 77486
rect 476805 77218 476847 77454
rect 477083 77218 477125 77454
rect 476805 77134 477125 77218
rect 476805 76898 476847 77134
rect 477083 76898 477125 77134
rect 476805 76866 477125 76898
rect 498874 77454 499194 77486
rect 498874 77218 498916 77454
rect 499152 77218 499194 77454
rect 498874 77134 499194 77218
rect 498874 76898 498916 77134
rect 499152 76898 499194 77134
rect 498874 76866 499194 76898
rect 504805 77454 505125 77486
rect 504805 77218 504847 77454
rect 505083 77218 505125 77454
rect 504805 77134 505125 77218
rect 504805 76898 504847 77134
rect 505083 76898 505125 77134
rect 504805 76866 505125 76898
rect 526874 77454 527194 77486
rect 526874 77218 526916 77454
rect 527152 77218 527194 77454
rect 526874 77134 527194 77218
rect 526874 76898 526916 77134
rect 527152 76898 527194 77134
rect 526874 76866 527194 76898
rect 532805 77454 533125 77486
rect 532805 77218 532847 77454
rect 533083 77218 533125 77454
rect 532805 77134 533125 77218
rect 532805 76898 532847 77134
rect 533083 76898 533125 77134
rect 532805 76866 533125 76898
rect 554874 77454 555194 77486
rect 554874 77218 554916 77454
rect 555152 77218 555194 77454
rect 554874 77134 555194 77218
rect 554874 76898 554916 77134
rect 555152 76898 555194 77134
rect 554874 76866 555194 76898
rect 560805 77454 561125 77486
rect 560805 77218 560847 77454
rect 561083 77218 561125 77454
rect 560805 77134 561125 77218
rect 560805 76898 560847 77134
rect 561083 76898 561125 77134
rect 560805 76866 561125 76898
rect -2006 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 -1386 53829
rect -2006 53509 -1386 53593
rect -2006 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 -1386 53509
rect -2006 26829 -1386 53273
rect 19910 53829 20230 53861
rect 19910 53593 19952 53829
rect 20188 53593 20230 53829
rect 19910 53509 20230 53593
rect 19910 53273 19952 53509
rect 20188 53273 20230 53509
rect 19910 53241 20230 53273
rect 25840 53829 26160 53861
rect 25840 53593 25882 53829
rect 26118 53593 26160 53829
rect 25840 53509 26160 53593
rect 25840 53273 25882 53509
rect 26118 53273 26160 53509
rect 25840 53241 26160 53273
rect 31771 53829 32091 53861
rect 31771 53593 31813 53829
rect 32049 53593 32091 53829
rect 31771 53509 32091 53593
rect 31771 53273 31813 53509
rect 32049 53273 32091 53509
rect 31771 53241 32091 53273
rect 47910 53829 48230 53861
rect 47910 53593 47952 53829
rect 48188 53593 48230 53829
rect 47910 53509 48230 53593
rect 47910 53273 47952 53509
rect 48188 53273 48230 53509
rect 47910 53241 48230 53273
rect 53840 53829 54160 53861
rect 53840 53593 53882 53829
rect 54118 53593 54160 53829
rect 53840 53509 54160 53593
rect 53840 53273 53882 53509
rect 54118 53273 54160 53509
rect 53840 53241 54160 53273
rect 59771 53829 60091 53861
rect 59771 53593 59813 53829
rect 60049 53593 60091 53829
rect 59771 53509 60091 53593
rect 59771 53273 59813 53509
rect 60049 53273 60091 53509
rect 59771 53241 60091 53273
rect 75910 53829 76230 53861
rect 75910 53593 75952 53829
rect 76188 53593 76230 53829
rect 75910 53509 76230 53593
rect 75910 53273 75952 53509
rect 76188 53273 76230 53509
rect 75910 53241 76230 53273
rect 81840 53829 82160 53861
rect 81840 53593 81882 53829
rect 82118 53593 82160 53829
rect 81840 53509 82160 53593
rect 81840 53273 81882 53509
rect 82118 53273 82160 53509
rect 81840 53241 82160 53273
rect 87771 53829 88091 53861
rect 87771 53593 87813 53829
rect 88049 53593 88091 53829
rect 87771 53509 88091 53593
rect 87771 53273 87813 53509
rect 88049 53273 88091 53509
rect 87771 53241 88091 53273
rect 103910 53829 104230 53861
rect 103910 53593 103952 53829
rect 104188 53593 104230 53829
rect 103910 53509 104230 53593
rect 103910 53273 103952 53509
rect 104188 53273 104230 53509
rect 103910 53241 104230 53273
rect 109840 53829 110160 53861
rect 109840 53593 109882 53829
rect 110118 53593 110160 53829
rect 109840 53509 110160 53593
rect 109840 53273 109882 53509
rect 110118 53273 110160 53509
rect 109840 53241 110160 53273
rect 115771 53829 116091 53861
rect 115771 53593 115813 53829
rect 116049 53593 116091 53829
rect 115771 53509 116091 53593
rect 115771 53273 115813 53509
rect 116049 53273 116091 53509
rect 115771 53241 116091 53273
rect 131910 53829 132230 53861
rect 131910 53593 131952 53829
rect 132188 53593 132230 53829
rect 131910 53509 132230 53593
rect 131910 53273 131952 53509
rect 132188 53273 132230 53509
rect 131910 53241 132230 53273
rect 137840 53829 138160 53861
rect 137840 53593 137882 53829
rect 138118 53593 138160 53829
rect 137840 53509 138160 53593
rect 137840 53273 137882 53509
rect 138118 53273 138160 53509
rect 137840 53241 138160 53273
rect 143771 53829 144091 53861
rect 143771 53593 143813 53829
rect 144049 53593 144091 53829
rect 143771 53509 144091 53593
rect 143771 53273 143813 53509
rect 144049 53273 144091 53509
rect 143771 53241 144091 53273
rect 159910 53829 160230 53861
rect 159910 53593 159952 53829
rect 160188 53593 160230 53829
rect 159910 53509 160230 53593
rect 159910 53273 159952 53509
rect 160188 53273 160230 53509
rect 159910 53241 160230 53273
rect 165840 53829 166160 53861
rect 165840 53593 165882 53829
rect 166118 53593 166160 53829
rect 165840 53509 166160 53593
rect 165840 53273 165882 53509
rect 166118 53273 166160 53509
rect 165840 53241 166160 53273
rect 171771 53829 172091 53861
rect 171771 53593 171813 53829
rect 172049 53593 172091 53829
rect 171771 53509 172091 53593
rect 171771 53273 171813 53509
rect 172049 53273 172091 53509
rect 171771 53241 172091 53273
rect 187910 53829 188230 53861
rect 187910 53593 187952 53829
rect 188188 53593 188230 53829
rect 187910 53509 188230 53593
rect 187910 53273 187952 53509
rect 188188 53273 188230 53509
rect 187910 53241 188230 53273
rect 193840 53829 194160 53861
rect 193840 53593 193882 53829
rect 194118 53593 194160 53829
rect 193840 53509 194160 53593
rect 193840 53273 193882 53509
rect 194118 53273 194160 53509
rect 193840 53241 194160 53273
rect 199771 53829 200091 53861
rect 199771 53593 199813 53829
rect 200049 53593 200091 53829
rect 199771 53509 200091 53593
rect 199771 53273 199813 53509
rect 200049 53273 200091 53509
rect 199771 53241 200091 53273
rect 215910 53829 216230 53861
rect 215910 53593 215952 53829
rect 216188 53593 216230 53829
rect 215910 53509 216230 53593
rect 215910 53273 215952 53509
rect 216188 53273 216230 53509
rect 215910 53241 216230 53273
rect 221840 53829 222160 53861
rect 221840 53593 221882 53829
rect 222118 53593 222160 53829
rect 221840 53509 222160 53593
rect 221840 53273 221882 53509
rect 222118 53273 222160 53509
rect 221840 53241 222160 53273
rect 227771 53829 228091 53861
rect 227771 53593 227813 53829
rect 228049 53593 228091 53829
rect 227771 53509 228091 53593
rect 227771 53273 227813 53509
rect 228049 53273 228091 53509
rect 227771 53241 228091 53273
rect 243910 53829 244230 53861
rect 243910 53593 243952 53829
rect 244188 53593 244230 53829
rect 243910 53509 244230 53593
rect 243910 53273 243952 53509
rect 244188 53273 244230 53509
rect 243910 53241 244230 53273
rect 249840 53829 250160 53861
rect 249840 53593 249882 53829
rect 250118 53593 250160 53829
rect 249840 53509 250160 53593
rect 249840 53273 249882 53509
rect 250118 53273 250160 53509
rect 249840 53241 250160 53273
rect 255771 53829 256091 53861
rect 255771 53593 255813 53829
rect 256049 53593 256091 53829
rect 255771 53509 256091 53593
rect 255771 53273 255813 53509
rect 256049 53273 256091 53509
rect 255771 53241 256091 53273
rect 271910 53829 272230 53861
rect 271910 53593 271952 53829
rect 272188 53593 272230 53829
rect 271910 53509 272230 53593
rect 271910 53273 271952 53509
rect 272188 53273 272230 53509
rect 271910 53241 272230 53273
rect 277840 53829 278160 53861
rect 277840 53593 277882 53829
rect 278118 53593 278160 53829
rect 277840 53509 278160 53593
rect 277840 53273 277882 53509
rect 278118 53273 278160 53509
rect 277840 53241 278160 53273
rect 283771 53829 284091 53861
rect 283771 53593 283813 53829
rect 284049 53593 284091 53829
rect 283771 53509 284091 53593
rect 283771 53273 283813 53509
rect 284049 53273 284091 53509
rect 283771 53241 284091 53273
rect 299910 53829 300230 53861
rect 299910 53593 299952 53829
rect 300188 53593 300230 53829
rect 299910 53509 300230 53593
rect 299910 53273 299952 53509
rect 300188 53273 300230 53509
rect 299910 53241 300230 53273
rect 305840 53829 306160 53861
rect 305840 53593 305882 53829
rect 306118 53593 306160 53829
rect 305840 53509 306160 53593
rect 305840 53273 305882 53509
rect 306118 53273 306160 53509
rect 305840 53241 306160 53273
rect 311771 53829 312091 53861
rect 311771 53593 311813 53829
rect 312049 53593 312091 53829
rect 311771 53509 312091 53593
rect 311771 53273 311813 53509
rect 312049 53273 312091 53509
rect 311771 53241 312091 53273
rect 327910 53829 328230 53861
rect 327910 53593 327952 53829
rect 328188 53593 328230 53829
rect 327910 53509 328230 53593
rect 327910 53273 327952 53509
rect 328188 53273 328230 53509
rect 327910 53241 328230 53273
rect 333840 53829 334160 53861
rect 333840 53593 333882 53829
rect 334118 53593 334160 53829
rect 333840 53509 334160 53593
rect 333840 53273 333882 53509
rect 334118 53273 334160 53509
rect 333840 53241 334160 53273
rect 339771 53829 340091 53861
rect 339771 53593 339813 53829
rect 340049 53593 340091 53829
rect 339771 53509 340091 53593
rect 339771 53273 339813 53509
rect 340049 53273 340091 53509
rect 339771 53241 340091 53273
rect 355910 53829 356230 53861
rect 355910 53593 355952 53829
rect 356188 53593 356230 53829
rect 355910 53509 356230 53593
rect 355910 53273 355952 53509
rect 356188 53273 356230 53509
rect 355910 53241 356230 53273
rect 361840 53829 362160 53861
rect 361840 53593 361882 53829
rect 362118 53593 362160 53829
rect 361840 53509 362160 53593
rect 361840 53273 361882 53509
rect 362118 53273 362160 53509
rect 361840 53241 362160 53273
rect 367771 53829 368091 53861
rect 367771 53593 367813 53829
rect 368049 53593 368091 53829
rect 367771 53509 368091 53593
rect 367771 53273 367813 53509
rect 368049 53273 368091 53509
rect 367771 53241 368091 53273
rect 383910 53829 384230 53861
rect 383910 53593 383952 53829
rect 384188 53593 384230 53829
rect 383910 53509 384230 53593
rect 383910 53273 383952 53509
rect 384188 53273 384230 53509
rect 383910 53241 384230 53273
rect 389840 53829 390160 53861
rect 389840 53593 389882 53829
rect 390118 53593 390160 53829
rect 389840 53509 390160 53593
rect 389840 53273 389882 53509
rect 390118 53273 390160 53509
rect 389840 53241 390160 53273
rect 395771 53829 396091 53861
rect 395771 53593 395813 53829
rect 396049 53593 396091 53829
rect 395771 53509 396091 53593
rect 395771 53273 395813 53509
rect 396049 53273 396091 53509
rect 395771 53241 396091 53273
rect 411910 53829 412230 53861
rect 411910 53593 411952 53829
rect 412188 53593 412230 53829
rect 411910 53509 412230 53593
rect 411910 53273 411952 53509
rect 412188 53273 412230 53509
rect 411910 53241 412230 53273
rect 417840 53829 418160 53861
rect 417840 53593 417882 53829
rect 418118 53593 418160 53829
rect 417840 53509 418160 53593
rect 417840 53273 417882 53509
rect 418118 53273 418160 53509
rect 417840 53241 418160 53273
rect 423771 53829 424091 53861
rect 423771 53593 423813 53829
rect 424049 53593 424091 53829
rect 423771 53509 424091 53593
rect 423771 53273 423813 53509
rect 424049 53273 424091 53509
rect 423771 53241 424091 53273
rect 439910 53829 440230 53861
rect 439910 53593 439952 53829
rect 440188 53593 440230 53829
rect 439910 53509 440230 53593
rect 439910 53273 439952 53509
rect 440188 53273 440230 53509
rect 439910 53241 440230 53273
rect 445840 53829 446160 53861
rect 445840 53593 445882 53829
rect 446118 53593 446160 53829
rect 445840 53509 446160 53593
rect 445840 53273 445882 53509
rect 446118 53273 446160 53509
rect 445840 53241 446160 53273
rect 451771 53829 452091 53861
rect 451771 53593 451813 53829
rect 452049 53593 452091 53829
rect 451771 53509 452091 53593
rect 451771 53273 451813 53509
rect 452049 53273 452091 53509
rect 451771 53241 452091 53273
rect 467910 53829 468230 53861
rect 467910 53593 467952 53829
rect 468188 53593 468230 53829
rect 467910 53509 468230 53593
rect 467910 53273 467952 53509
rect 468188 53273 468230 53509
rect 467910 53241 468230 53273
rect 473840 53829 474160 53861
rect 473840 53593 473882 53829
rect 474118 53593 474160 53829
rect 473840 53509 474160 53593
rect 473840 53273 473882 53509
rect 474118 53273 474160 53509
rect 473840 53241 474160 53273
rect 479771 53829 480091 53861
rect 479771 53593 479813 53829
rect 480049 53593 480091 53829
rect 479771 53509 480091 53593
rect 479771 53273 479813 53509
rect 480049 53273 480091 53509
rect 479771 53241 480091 53273
rect 495910 53829 496230 53861
rect 495910 53593 495952 53829
rect 496188 53593 496230 53829
rect 495910 53509 496230 53593
rect 495910 53273 495952 53509
rect 496188 53273 496230 53509
rect 495910 53241 496230 53273
rect 501840 53829 502160 53861
rect 501840 53593 501882 53829
rect 502118 53593 502160 53829
rect 501840 53509 502160 53593
rect 501840 53273 501882 53509
rect 502118 53273 502160 53509
rect 501840 53241 502160 53273
rect 507771 53829 508091 53861
rect 507771 53593 507813 53829
rect 508049 53593 508091 53829
rect 507771 53509 508091 53593
rect 507771 53273 507813 53509
rect 508049 53273 508091 53509
rect 507771 53241 508091 53273
rect 523910 53829 524230 53861
rect 523910 53593 523952 53829
rect 524188 53593 524230 53829
rect 523910 53509 524230 53593
rect 523910 53273 523952 53509
rect 524188 53273 524230 53509
rect 523910 53241 524230 53273
rect 529840 53829 530160 53861
rect 529840 53593 529882 53829
rect 530118 53593 530160 53829
rect 529840 53509 530160 53593
rect 529840 53273 529882 53509
rect 530118 53273 530160 53509
rect 529840 53241 530160 53273
rect 535771 53829 536091 53861
rect 535771 53593 535813 53829
rect 536049 53593 536091 53829
rect 535771 53509 536091 53593
rect 535771 53273 535813 53509
rect 536049 53273 536091 53509
rect 535771 53241 536091 53273
rect 551910 53829 552230 53861
rect 551910 53593 551952 53829
rect 552188 53593 552230 53829
rect 551910 53509 552230 53593
rect 551910 53273 551952 53509
rect 552188 53273 552230 53509
rect 551910 53241 552230 53273
rect 557840 53829 558160 53861
rect 557840 53593 557882 53829
rect 558118 53593 558160 53829
rect 557840 53509 558160 53593
rect 557840 53273 557882 53509
rect 558118 53273 558160 53509
rect 557840 53241 558160 53273
rect 563771 53829 564091 53861
rect 563771 53593 563813 53829
rect 564049 53593 564091 53829
rect 563771 53509 564091 53593
rect 563771 53273 563813 53509
rect 564049 53273 564091 53509
rect 563771 53241 564091 53273
rect 573494 53829 574114 80273
rect 573494 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 574114 53829
rect 573494 53509 574114 53593
rect 573494 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 574114 53509
rect 22874 50454 23194 50486
rect 22874 50218 22916 50454
rect 23152 50218 23194 50454
rect 22874 50134 23194 50218
rect 22874 49898 22916 50134
rect 23152 49898 23194 50134
rect 22874 49866 23194 49898
rect 28805 50454 29125 50486
rect 28805 50218 28847 50454
rect 29083 50218 29125 50454
rect 28805 50134 29125 50218
rect 28805 49898 28847 50134
rect 29083 49898 29125 50134
rect 28805 49866 29125 49898
rect 50874 50454 51194 50486
rect 50874 50218 50916 50454
rect 51152 50218 51194 50454
rect 50874 50134 51194 50218
rect 50874 49898 50916 50134
rect 51152 49898 51194 50134
rect 50874 49866 51194 49898
rect 56805 50454 57125 50486
rect 56805 50218 56847 50454
rect 57083 50218 57125 50454
rect 56805 50134 57125 50218
rect 56805 49898 56847 50134
rect 57083 49898 57125 50134
rect 56805 49866 57125 49898
rect 78874 50454 79194 50486
rect 78874 50218 78916 50454
rect 79152 50218 79194 50454
rect 78874 50134 79194 50218
rect 78874 49898 78916 50134
rect 79152 49898 79194 50134
rect 78874 49866 79194 49898
rect 84805 50454 85125 50486
rect 84805 50218 84847 50454
rect 85083 50218 85125 50454
rect 84805 50134 85125 50218
rect 84805 49898 84847 50134
rect 85083 49898 85125 50134
rect 84805 49866 85125 49898
rect 106874 50454 107194 50486
rect 106874 50218 106916 50454
rect 107152 50218 107194 50454
rect 106874 50134 107194 50218
rect 106874 49898 106916 50134
rect 107152 49898 107194 50134
rect 106874 49866 107194 49898
rect 112805 50454 113125 50486
rect 112805 50218 112847 50454
rect 113083 50218 113125 50454
rect 112805 50134 113125 50218
rect 112805 49898 112847 50134
rect 113083 49898 113125 50134
rect 112805 49866 113125 49898
rect 134874 50454 135194 50486
rect 134874 50218 134916 50454
rect 135152 50218 135194 50454
rect 134874 50134 135194 50218
rect 134874 49898 134916 50134
rect 135152 49898 135194 50134
rect 134874 49866 135194 49898
rect 140805 50454 141125 50486
rect 140805 50218 140847 50454
rect 141083 50218 141125 50454
rect 140805 50134 141125 50218
rect 140805 49898 140847 50134
rect 141083 49898 141125 50134
rect 140805 49866 141125 49898
rect 162874 50454 163194 50486
rect 162874 50218 162916 50454
rect 163152 50218 163194 50454
rect 162874 50134 163194 50218
rect 162874 49898 162916 50134
rect 163152 49898 163194 50134
rect 162874 49866 163194 49898
rect 168805 50454 169125 50486
rect 168805 50218 168847 50454
rect 169083 50218 169125 50454
rect 168805 50134 169125 50218
rect 168805 49898 168847 50134
rect 169083 49898 169125 50134
rect 168805 49866 169125 49898
rect 190874 50454 191194 50486
rect 190874 50218 190916 50454
rect 191152 50218 191194 50454
rect 190874 50134 191194 50218
rect 190874 49898 190916 50134
rect 191152 49898 191194 50134
rect 190874 49866 191194 49898
rect 196805 50454 197125 50486
rect 196805 50218 196847 50454
rect 197083 50218 197125 50454
rect 196805 50134 197125 50218
rect 196805 49898 196847 50134
rect 197083 49898 197125 50134
rect 196805 49866 197125 49898
rect 218874 50454 219194 50486
rect 218874 50218 218916 50454
rect 219152 50218 219194 50454
rect 218874 50134 219194 50218
rect 218874 49898 218916 50134
rect 219152 49898 219194 50134
rect 218874 49866 219194 49898
rect 224805 50454 225125 50486
rect 224805 50218 224847 50454
rect 225083 50218 225125 50454
rect 224805 50134 225125 50218
rect 224805 49898 224847 50134
rect 225083 49898 225125 50134
rect 224805 49866 225125 49898
rect 246874 50454 247194 50486
rect 246874 50218 246916 50454
rect 247152 50218 247194 50454
rect 246874 50134 247194 50218
rect 246874 49898 246916 50134
rect 247152 49898 247194 50134
rect 246874 49866 247194 49898
rect 252805 50454 253125 50486
rect 252805 50218 252847 50454
rect 253083 50218 253125 50454
rect 252805 50134 253125 50218
rect 252805 49898 252847 50134
rect 253083 49898 253125 50134
rect 252805 49866 253125 49898
rect 274874 50454 275194 50486
rect 274874 50218 274916 50454
rect 275152 50218 275194 50454
rect 274874 50134 275194 50218
rect 274874 49898 274916 50134
rect 275152 49898 275194 50134
rect 274874 49866 275194 49898
rect 280805 50454 281125 50486
rect 280805 50218 280847 50454
rect 281083 50218 281125 50454
rect 280805 50134 281125 50218
rect 280805 49898 280847 50134
rect 281083 49898 281125 50134
rect 280805 49866 281125 49898
rect 302874 50454 303194 50486
rect 302874 50218 302916 50454
rect 303152 50218 303194 50454
rect 302874 50134 303194 50218
rect 302874 49898 302916 50134
rect 303152 49898 303194 50134
rect 302874 49866 303194 49898
rect 308805 50454 309125 50486
rect 308805 50218 308847 50454
rect 309083 50218 309125 50454
rect 308805 50134 309125 50218
rect 308805 49898 308847 50134
rect 309083 49898 309125 50134
rect 308805 49866 309125 49898
rect 330874 50454 331194 50486
rect 330874 50218 330916 50454
rect 331152 50218 331194 50454
rect 330874 50134 331194 50218
rect 330874 49898 330916 50134
rect 331152 49898 331194 50134
rect 330874 49866 331194 49898
rect 336805 50454 337125 50486
rect 336805 50218 336847 50454
rect 337083 50218 337125 50454
rect 336805 50134 337125 50218
rect 336805 49898 336847 50134
rect 337083 49898 337125 50134
rect 336805 49866 337125 49898
rect 358874 50454 359194 50486
rect 358874 50218 358916 50454
rect 359152 50218 359194 50454
rect 358874 50134 359194 50218
rect 358874 49898 358916 50134
rect 359152 49898 359194 50134
rect 358874 49866 359194 49898
rect 364805 50454 365125 50486
rect 364805 50218 364847 50454
rect 365083 50218 365125 50454
rect 364805 50134 365125 50218
rect 364805 49898 364847 50134
rect 365083 49898 365125 50134
rect 364805 49866 365125 49898
rect 386874 50454 387194 50486
rect 386874 50218 386916 50454
rect 387152 50218 387194 50454
rect 386874 50134 387194 50218
rect 386874 49898 386916 50134
rect 387152 49898 387194 50134
rect 386874 49866 387194 49898
rect 392805 50454 393125 50486
rect 392805 50218 392847 50454
rect 393083 50218 393125 50454
rect 392805 50134 393125 50218
rect 392805 49898 392847 50134
rect 393083 49898 393125 50134
rect 392805 49866 393125 49898
rect 414874 50454 415194 50486
rect 414874 50218 414916 50454
rect 415152 50218 415194 50454
rect 414874 50134 415194 50218
rect 414874 49898 414916 50134
rect 415152 49898 415194 50134
rect 414874 49866 415194 49898
rect 420805 50454 421125 50486
rect 420805 50218 420847 50454
rect 421083 50218 421125 50454
rect 420805 50134 421125 50218
rect 420805 49898 420847 50134
rect 421083 49898 421125 50134
rect 420805 49866 421125 49898
rect 442874 50454 443194 50486
rect 442874 50218 442916 50454
rect 443152 50218 443194 50454
rect 442874 50134 443194 50218
rect 442874 49898 442916 50134
rect 443152 49898 443194 50134
rect 442874 49866 443194 49898
rect 448805 50454 449125 50486
rect 448805 50218 448847 50454
rect 449083 50218 449125 50454
rect 448805 50134 449125 50218
rect 448805 49898 448847 50134
rect 449083 49898 449125 50134
rect 448805 49866 449125 49898
rect 470874 50454 471194 50486
rect 470874 50218 470916 50454
rect 471152 50218 471194 50454
rect 470874 50134 471194 50218
rect 470874 49898 470916 50134
rect 471152 49898 471194 50134
rect 470874 49866 471194 49898
rect 476805 50454 477125 50486
rect 476805 50218 476847 50454
rect 477083 50218 477125 50454
rect 476805 50134 477125 50218
rect 476805 49898 476847 50134
rect 477083 49898 477125 50134
rect 476805 49866 477125 49898
rect 498874 50454 499194 50486
rect 498874 50218 498916 50454
rect 499152 50218 499194 50454
rect 498874 50134 499194 50218
rect 498874 49898 498916 50134
rect 499152 49898 499194 50134
rect 498874 49866 499194 49898
rect 504805 50454 505125 50486
rect 504805 50218 504847 50454
rect 505083 50218 505125 50454
rect 504805 50134 505125 50218
rect 504805 49898 504847 50134
rect 505083 49898 505125 50134
rect 504805 49866 505125 49898
rect 526874 50454 527194 50486
rect 526874 50218 526916 50454
rect 527152 50218 527194 50454
rect 526874 50134 527194 50218
rect 526874 49898 526916 50134
rect 527152 49898 527194 50134
rect 526874 49866 527194 49898
rect 532805 50454 533125 50486
rect 532805 50218 532847 50454
rect 533083 50218 533125 50454
rect 532805 50134 533125 50218
rect 532805 49898 532847 50134
rect 533083 49898 533125 50134
rect 532805 49866 533125 49898
rect 554874 50454 555194 50486
rect 554874 50218 554916 50454
rect 555152 50218 555194 50454
rect 554874 50134 555194 50218
rect 554874 49898 554916 50134
rect 555152 49898 555194 50134
rect 554874 49866 555194 49898
rect 560805 50454 561125 50486
rect 560805 50218 560847 50454
rect 561083 50218 561125 50454
rect 560805 50134 561125 50218
rect 560805 49898 560847 50134
rect 561083 49898 561125 50134
rect 560805 49866 561125 49898
rect -2006 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 -1386 26829
rect -2006 26509 -1386 26593
rect -2006 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 -1386 26509
rect -2006 -346 -1386 26273
rect 24242 26829 24562 26861
rect 24242 26593 24284 26829
rect 24520 26593 24562 26829
rect 24242 26509 24562 26593
rect 24242 26273 24284 26509
rect 24520 26273 24562 26509
rect 24242 26241 24562 26273
rect 38840 26829 39160 26861
rect 38840 26593 38882 26829
rect 39118 26593 39160 26829
rect 38840 26509 39160 26593
rect 38840 26273 38882 26509
rect 39118 26273 39160 26509
rect 38840 26241 39160 26273
rect 53437 26829 53757 26861
rect 53437 26593 53479 26829
rect 53715 26593 53757 26829
rect 53437 26509 53757 26593
rect 53437 26273 53479 26509
rect 53715 26273 53757 26509
rect 53437 26241 53757 26273
rect 31542 23454 31862 23486
rect 31542 23218 31584 23454
rect 31820 23218 31862 23454
rect 31542 23134 31862 23218
rect 31542 22898 31584 23134
rect 31820 22898 31862 23134
rect 31542 22866 31862 22898
rect 46139 23454 46459 23486
rect 46139 23218 46181 23454
rect 46417 23218 46459 23454
rect 46139 23134 46459 23218
rect 46139 22898 46181 23134
rect 46417 22898 46459 23134
rect 46139 22866 46459 22898
rect 65994 23454 66614 41000
rect 75910 26829 76230 26861
rect 75910 26593 75952 26829
rect 76188 26593 76230 26829
rect 75910 26509 76230 26593
rect 75910 26273 75952 26509
rect 76188 26273 76230 26509
rect 75910 26241 76230 26273
rect 81840 26829 82160 26861
rect 81840 26593 81882 26829
rect 82118 26593 82160 26829
rect 81840 26509 82160 26593
rect 81840 26273 81882 26509
rect 82118 26273 82160 26509
rect 81840 26241 82160 26273
rect 87771 26829 88091 26861
rect 87771 26593 87813 26829
rect 88049 26593 88091 26829
rect 87771 26509 88091 26593
rect 87771 26273 87813 26509
rect 88049 26273 88091 26509
rect 87771 26241 88091 26273
rect 103910 26829 104230 26861
rect 103910 26593 103952 26829
rect 104188 26593 104230 26829
rect 103910 26509 104230 26593
rect 103910 26273 103952 26509
rect 104188 26273 104230 26509
rect 103910 26241 104230 26273
rect 109840 26829 110160 26861
rect 109840 26593 109882 26829
rect 110118 26593 110160 26829
rect 109840 26509 110160 26593
rect 109840 26273 109882 26509
rect 110118 26273 110160 26509
rect 109840 26241 110160 26273
rect 115771 26829 116091 26861
rect 115771 26593 115813 26829
rect 116049 26593 116091 26829
rect 115771 26509 116091 26593
rect 115771 26273 115813 26509
rect 116049 26273 116091 26509
rect 115771 26241 116091 26273
rect 131910 26829 132230 26861
rect 131910 26593 131952 26829
rect 132188 26593 132230 26829
rect 131910 26509 132230 26593
rect 131910 26273 131952 26509
rect 132188 26273 132230 26509
rect 131910 26241 132230 26273
rect 137840 26829 138160 26861
rect 137840 26593 137882 26829
rect 138118 26593 138160 26829
rect 137840 26509 138160 26593
rect 137840 26273 137882 26509
rect 138118 26273 138160 26509
rect 137840 26241 138160 26273
rect 143771 26829 144091 26861
rect 143771 26593 143813 26829
rect 144049 26593 144091 26829
rect 143771 26509 144091 26593
rect 143771 26273 143813 26509
rect 144049 26273 144091 26509
rect 143771 26241 144091 26273
rect 159910 26829 160230 26861
rect 159910 26593 159952 26829
rect 160188 26593 160230 26829
rect 159910 26509 160230 26593
rect 159910 26273 159952 26509
rect 160188 26273 160230 26509
rect 159910 26241 160230 26273
rect 165840 26829 166160 26861
rect 165840 26593 165882 26829
rect 166118 26593 166160 26829
rect 165840 26509 166160 26593
rect 165840 26273 165882 26509
rect 166118 26273 166160 26509
rect 165840 26241 166160 26273
rect 171771 26829 172091 26861
rect 171771 26593 171813 26829
rect 172049 26593 172091 26829
rect 171771 26509 172091 26593
rect 171771 26273 171813 26509
rect 172049 26273 172091 26509
rect 171771 26241 172091 26273
rect 187910 26829 188230 26861
rect 187910 26593 187952 26829
rect 188188 26593 188230 26829
rect 187910 26509 188230 26593
rect 187910 26273 187952 26509
rect 188188 26273 188230 26509
rect 187910 26241 188230 26273
rect 193840 26829 194160 26861
rect 193840 26593 193882 26829
rect 194118 26593 194160 26829
rect 193840 26509 194160 26593
rect 193840 26273 193882 26509
rect 194118 26273 194160 26509
rect 193840 26241 194160 26273
rect 199771 26829 200091 26861
rect 199771 26593 199813 26829
rect 200049 26593 200091 26829
rect 199771 26509 200091 26593
rect 199771 26273 199813 26509
rect 200049 26273 200091 26509
rect 199771 26241 200091 26273
rect 215910 26829 216230 26861
rect 215910 26593 215952 26829
rect 216188 26593 216230 26829
rect 215910 26509 216230 26593
rect 215910 26273 215952 26509
rect 216188 26273 216230 26509
rect 215910 26241 216230 26273
rect 221840 26829 222160 26861
rect 221840 26593 221882 26829
rect 222118 26593 222160 26829
rect 221840 26509 222160 26593
rect 221840 26273 221882 26509
rect 222118 26273 222160 26509
rect 221840 26241 222160 26273
rect 227771 26829 228091 26861
rect 227771 26593 227813 26829
rect 228049 26593 228091 26829
rect 227771 26509 228091 26593
rect 227771 26273 227813 26509
rect 228049 26273 228091 26509
rect 227771 26241 228091 26273
rect 243910 26829 244230 26861
rect 243910 26593 243952 26829
rect 244188 26593 244230 26829
rect 243910 26509 244230 26593
rect 243910 26273 243952 26509
rect 244188 26273 244230 26509
rect 243910 26241 244230 26273
rect 249840 26829 250160 26861
rect 249840 26593 249882 26829
rect 250118 26593 250160 26829
rect 249840 26509 250160 26593
rect 249840 26273 249882 26509
rect 250118 26273 250160 26509
rect 249840 26241 250160 26273
rect 255771 26829 256091 26861
rect 255771 26593 255813 26829
rect 256049 26593 256091 26829
rect 255771 26509 256091 26593
rect 255771 26273 255813 26509
rect 256049 26273 256091 26509
rect 255771 26241 256091 26273
rect 271910 26829 272230 26861
rect 271910 26593 271952 26829
rect 272188 26593 272230 26829
rect 271910 26509 272230 26593
rect 271910 26273 271952 26509
rect 272188 26273 272230 26509
rect 271910 26241 272230 26273
rect 277840 26829 278160 26861
rect 277840 26593 277882 26829
rect 278118 26593 278160 26829
rect 277840 26509 278160 26593
rect 277840 26273 277882 26509
rect 278118 26273 278160 26509
rect 277840 26241 278160 26273
rect 283771 26829 284091 26861
rect 283771 26593 283813 26829
rect 284049 26593 284091 26829
rect 283771 26509 284091 26593
rect 283771 26273 283813 26509
rect 284049 26273 284091 26509
rect 283771 26241 284091 26273
rect 299910 26829 300230 26861
rect 299910 26593 299952 26829
rect 300188 26593 300230 26829
rect 299910 26509 300230 26593
rect 299910 26273 299952 26509
rect 300188 26273 300230 26509
rect 299910 26241 300230 26273
rect 305840 26829 306160 26861
rect 305840 26593 305882 26829
rect 306118 26593 306160 26829
rect 305840 26509 306160 26593
rect 305840 26273 305882 26509
rect 306118 26273 306160 26509
rect 305840 26241 306160 26273
rect 311771 26829 312091 26861
rect 311771 26593 311813 26829
rect 312049 26593 312091 26829
rect 311771 26509 312091 26593
rect 311771 26273 311813 26509
rect 312049 26273 312091 26509
rect 311771 26241 312091 26273
rect 327910 26829 328230 26861
rect 327910 26593 327952 26829
rect 328188 26593 328230 26829
rect 327910 26509 328230 26593
rect 327910 26273 327952 26509
rect 328188 26273 328230 26509
rect 327910 26241 328230 26273
rect 333840 26829 334160 26861
rect 333840 26593 333882 26829
rect 334118 26593 334160 26829
rect 333840 26509 334160 26593
rect 333840 26273 333882 26509
rect 334118 26273 334160 26509
rect 333840 26241 334160 26273
rect 339771 26829 340091 26861
rect 339771 26593 339813 26829
rect 340049 26593 340091 26829
rect 339771 26509 340091 26593
rect 339771 26273 339813 26509
rect 340049 26273 340091 26509
rect 339771 26241 340091 26273
rect 355910 26829 356230 26861
rect 355910 26593 355952 26829
rect 356188 26593 356230 26829
rect 355910 26509 356230 26593
rect 355910 26273 355952 26509
rect 356188 26273 356230 26509
rect 355910 26241 356230 26273
rect 361840 26829 362160 26861
rect 361840 26593 361882 26829
rect 362118 26593 362160 26829
rect 361840 26509 362160 26593
rect 361840 26273 361882 26509
rect 362118 26273 362160 26509
rect 361840 26241 362160 26273
rect 367771 26829 368091 26861
rect 367771 26593 367813 26829
rect 368049 26593 368091 26829
rect 367771 26509 368091 26593
rect 367771 26273 367813 26509
rect 368049 26273 368091 26509
rect 367771 26241 368091 26273
rect 383910 26829 384230 26861
rect 383910 26593 383952 26829
rect 384188 26593 384230 26829
rect 383910 26509 384230 26593
rect 383910 26273 383952 26509
rect 384188 26273 384230 26509
rect 383910 26241 384230 26273
rect 389840 26829 390160 26861
rect 389840 26593 389882 26829
rect 390118 26593 390160 26829
rect 389840 26509 390160 26593
rect 389840 26273 389882 26509
rect 390118 26273 390160 26509
rect 389840 26241 390160 26273
rect 395771 26829 396091 26861
rect 395771 26593 395813 26829
rect 396049 26593 396091 26829
rect 395771 26509 396091 26593
rect 395771 26273 395813 26509
rect 396049 26273 396091 26509
rect 395771 26241 396091 26273
rect 411910 26829 412230 26861
rect 411910 26593 411952 26829
rect 412188 26593 412230 26829
rect 411910 26509 412230 26593
rect 411910 26273 411952 26509
rect 412188 26273 412230 26509
rect 411910 26241 412230 26273
rect 417840 26829 418160 26861
rect 417840 26593 417882 26829
rect 418118 26593 418160 26829
rect 417840 26509 418160 26593
rect 417840 26273 417882 26509
rect 418118 26273 418160 26509
rect 417840 26241 418160 26273
rect 423771 26829 424091 26861
rect 423771 26593 423813 26829
rect 424049 26593 424091 26829
rect 423771 26509 424091 26593
rect 423771 26273 423813 26509
rect 424049 26273 424091 26509
rect 423771 26241 424091 26273
rect 439910 26829 440230 26861
rect 439910 26593 439952 26829
rect 440188 26593 440230 26829
rect 439910 26509 440230 26593
rect 439910 26273 439952 26509
rect 440188 26273 440230 26509
rect 439910 26241 440230 26273
rect 445840 26829 446160 26861
rect 445840 26593 445882 26829
rect 446118 26593 446160 26829
rect 445840 26509 446160 26593
rect 445840 26273 445882 26509
rect 446118 26273 446160 26509
rect 445840 26241 446160 26273
rect 451771 26829 452091 26861
rect 451771 26593 451813 26829
rect 452049 26593 452091 26829
rect 451771 26509 452091 26593
rect 451771 26273 451813 26509
rect 452049 26273 452091 26509
rect 451771 26241 452091 26273
rect 467910 26829 468230 26861
rect 467910 26593 467952 26829
rect 468188 26593 468230 26829
rect 467910 26509 468230 26593
rect 467910 26273 467952 26509
rect 468188 26273 468230 26509
rect 467910 26241 468230 26273
rect 473840 26829 474160 26861
rect 473840 26593 473882 26829
rect 474118 26593 474160 26829
rect 473840 26509 474160 26593
rect 473840 26273 473882 26509
rect 474118 26273 474160 26509
rect 473840 26241 474160 26273
rect 479771 26829 480091 26861
rect 479771 26593 479813 26829
rect 480049 26593 480091 26829
rect 479771 26509 480091 26593
rect 479771 26273 479813 26509
rect 480049 26273 480091 26509
rect 479771 26241 480091 26273
rect 495910 26829 496230 26861
rect 495910 26593 495952 26829
rect 496188 26593 496230 26829
rect 495910 26509 496230 26593
rect 495910 26273 495952 26509
rect 496188 26273 496230 26509
rect 495910 26241 496230 26273
rect 501840 26829 502160 26861
rect 501840 26593 501882 26829
rect 502118 26593 502160 26829
rect 501840 26509 502160 26593
rect 501840 26273 501882 26509
rect 502118 26273 502160 26509
rect 501840 26241 502160 26273
rect 507771 26829 508091 26861
rect 507771 26593 507813 26829
rect 508049 26593 508091 26829
rect 507771 26509 508091 26593
rect 507771 26273 507813 26509
rect 508049 26273 508091 26509
rect 507771 26241 508091 26273
rect 523910 26829 524230 26861
rect 523910 26593 523952 26829
rect 524188 26593 524230 26829
rect 523910 26509 524230 26593
rect 523910 26273 523952 26509
rect 524188 26273 524230 26509
rect 523910 26241 524230 26273
rect 529840 26829 530160 26861
rect 529840 26593 529882 26829
rect 530118 26593 530160 26829
rect 529840 26509 530160 26593
rect 529840 26273 529882 26509
rect 530118 26273 530160 26509
rect 529840 26241 530160 26273
rect 535771 26829 536091 26861
rect 535771 26593 535813 26829
rect 536049 26593 536091 26829
rect 535771 26509 536091 26593
rect 535771 26273 535813 26509
rect 536049 26273 536091 26509
rect 535771 26241 536091 26273
rect 551910 26829 552230 26861
rect 551910 26593 551952 26829
rect 552188 26593 552230 26829
rect 551910 26509 552230 26593
rect 551910 26273 551952 26509
rect 552188 26273 552230 26509
rect 551910 26241 552230 26273
rect 557840 26829 558160 26861
rect 557840 26593 557882 26829
rect 558118 26593 558160 26829
rect 557840 26509 558160 26593
rect 557840 26273 557882 26509
rect 558118 26273 558160 26509
rect 557840 26241 558160 26273
rect 563771 26829 564091 26861
rect 563771 26593 563813 26829
rect 564049 26593 564091 26829
rect 563771 26509 564091 26593
rect 563771 26273 563813 26509
rect 564049 26273 564091 26509
rect 563771 26241 564091 26273
rect 573494 26829 574114 53273
rect 573494 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 574114 26829
rect 573494 26509 574114 26593
rect 573494 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 574114 26509
rect 65994 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 66614 23454
rect 65994 23134 66614 23218
rect 65994 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 66614 23134
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 65994 -1306 66614 22898
rect 78874 23454 79194 23486
rect 78874 23218 78916 23454
rect 79152 23218 79194 23454
rect 78874 23134 79194 23218
rect 78874 22898 78916 23134
rect 79152 22898 79194 23134
rect 78874 22866 79194 22898
rect 84805 23454 85125 23486
rect 84805 23218 84847 23454
rect 85083 23218 85125 23454
rect 84805 23134 85125 23218
rect 84805 22898 84847 23134
rect 85083 22898 85125 23134
rect 84805 22866 85125 22898
rect 106874 23454 107194 23486
rect 106874 23218 106916 23454
rect 107152 23218 107194 23454
rect 106874 23134 107194 23218
rect 106874 22898 106916 23134
rect 107152 22898 107194 23134
rect 106874 22866 107194 22898
rect 112805 23454 113125 23486
rect 112805 23218 112847 23454
rect 113083 23218 113125 23454
rect 112805 23134 113125 23218
rect 112805 22898 112847 23134
rect 113083 22898 113125 23134
rect 112805 22866 113125 22898
rect 134874 23454 135194 23486
rect 134874 23218 134916 23454
rect 135152 23218 135194 23454
rect 134874 23134 135194 23218
rect 134874 22898 134916 23134
rect 135152 22898 135194 23134
rect 134874 22866 135194 22898
rect 140805 23454 141125 23486
rect 140805 23218 140847 23454
rect 141083 23218 141125 23454
rect 140805 23134 141125 23218
rect 140805 22898 140847 23134
rect 141083 22898 141125 23134
rect 140805 22866 141125 22898
rect 162874 23454 163194 23486
rect 162874 23218 162916 23454
rect 163152 23218 163194 23454
rect 162874 23134 163194 23218
rect 162874 22898 162916 23134
rect 163152 22898 163194 23134
rect 162874 22866 163194 22898
rect 168805 23454 169125 23486
rect 168805 23218 168847 23454
rect 169083 23218 169125 23454
rect 168805 23134 169125 23218
rect 168805 22898 168847 23134
rect 169083 22898 169125 23134
rect 168805 22866 169125 22898
rect 190874 23454 191194 23486
rect 190874 23218 190916 23454
rect 191152 23218 191194 23454
rect 190874 23134 191194 23218
rect 190874 22898 190916 23134
rect 191152 22898 191194 23134
rect 190874 22866 191194 22898
rect 196805 23454 197125 23486
rect 196805 23218 196847 23454
rect 197083 23218 197125 23454
rect 196805 23134 197125 23218
rect 196805 22898 196847 23134
rect 197083 22898 197125 23134
rect 196805 22866 197125 22898
rect 218874 23454 219194 23486
rect 218874 23218 218916 23454
rect 219152 23218 219194 23454
rect 218874 23134 219194 23218
rect 218874 22898 218916 23134
rect 219152 22898 219194 23134
rect 218874 22866 219194 22898
rect 224805 23454 225125 23486
rect 224805 23218 224847 23454
rect 225083 23218 225125 23454
rect 224805 23134 225125 23218
rect 224805 22898 224847 23134
rect 225083 22898 225125 23134
rect 224805 22866 225125 22898
rect 246874 23454 247194 23486
rect 246874 23218 246916 23454
rect 247152 23218 247194 23454
rect 246874 23134 247194 23218
rect 246874 22898 246916 23134
rect 247152 22898 247194 23134
rect 246874 22866 247194 22898
rect 252805 23454 253125 23486
rect 252805 23218 252847 23454
rect 253083 23218 253125 23454
rect 252805 23134 253125 23218
rect 252805 22898 252847 23134
rect 253083 22898 253125 23134
rect 252805 22866 253125 22898
rect 274874 23454 275194 23486
rect 274874 23218 274916 23454
rect 275152 23218 275194 23454
rect 274874 23134 275194 23218
rect 274874 22898 274916 23134
rect 275152 22898 275194 23134
rect 274874 22866 275194 22898
rect 280805 23454 281125 23486
rect 280805 23218 280847 23454
rect 281083 23218 281125 23454
rect 280805 23134 281125 23218
rect 280805 22898 280847 23134
rect 281083 22898 281125 23134
rect 280805 22866 281125 22898
rect 302874 23454 303194 23486
rect 302874 23218 302916 23454
rect 303152 23218 303194 23454
rect 302874 23134 303194 23218
rect 302874 22898 302916 23134
rect 303152 22898 303194 23134
rect 302874 22866 303194 22898
rect 308805 23454 309125 23486
rect 308805 23218 308847 23454
rect 309083 23218 309125 23454
rect 308805 23134 309125 23218
rect 308805 22898 308847 23134
rect 309083 22898 309125 23134
rect 308805 22866 309125 22898
rect 330874 23454 331194 23486
rect 330874 23218 330916 23454
rect 331152 23218 331194 23454
rect 330874 23134 331194 23218
rect 330874 22898 330916 23134
rect 331152 22898 331194 23134
rect 330874 22866 331194 22898
rect 336805 23454 337125 23486
rect 336805 23218 336847 23454
rect 337083 23218 337125 23454
rect 336805 23134 337125 23218
rect 336805 22898 336847 23134
rect 337083 22898 337125 23134
rect 336805 22866 337125 22898
rect 358874 23454 359194 23486
rect 358874 23218 358916 23454
rect 359152 23218 359194 23454
rect 358874 23134 359194 23218
rect 358874 22898 358916 23134
rect 359152 22898 359194 23134
rect 358874 22866 359194 22898
rect 364805 23454 365125 23486
rect 364805 23218 364847 23454
rect 365083 23218 365125 23454
rect 364805 23134 365125 23218
rect 364805 22898 364847 23134
rect 365083 22898 365125 23134
rect 364805 22866 365125 22898
rect 386874 23454 387194 23486
rect 386874 23218 386916 23454
rect 387152 23218 387194 23454
rect 386874 23134 387194 23218
rect 386874 22898 386916 23134
rect 387152 22898 387194 23134
rect 386874 22866 387194 22898
rect 392805 23454 393125 23486
rect 392805 23218 392847 23454
rect 393083 23218 393125 23454
rect 392805 23134 393125 23218
rect 392805 22898 392847 23134
rect 393083 22898 393125 23134
rect 392805 22866 393125 22898
rect 414874 23454 415194 23486
rect 414874 23218 414916 23454
rect 415152 23218 415194 23454
rect 414874 23134 415194 23218
rect 414874 22898 414916 23134
rect 415152 22898 415194 23134
rect 414874 22866 415194 22898
rect 420805 23454 421125 23486
rect 420805 23218 420847 23454
rect 421083 23218 421125 23454
rect 420805 23134 421125 23218
rect 420805 22898 420847 23134
rect 421083 22898 421125 23134
rect 420805 22866 421125 22898
rect 442874 23454 443194 23486
rect 442874 23218 442916 23454
rect 443152 23218 443194 23454
rect 442874 23134 443194 23218
rect 442874 22898 442916 23134
rect 443152 22898 443194 23134
rect 442874 22866 443194 22898
rect 448805 23454 449125 23486
rect 448805 23218 448847 23454
rect 449083 23218 449125 23454
rect 448805 23134 449125 23218
rect 448805 22898 448847 23134
rect 449083 22898 449125 23134
rect 448805 22866 449125 22898
rect 470874 23454 471194 23486
rect 470874 23218 470916 23454
rect 471152 23218 471194 23454
rect 470874 23134 471194 23218
rect 470874 22898 470916 23134
rect 471152 22898 471194 23134
rect 470874 22866 471194 22898
rect 476805 23454 477125 23486
rect 476805 23218 476847 23454
rect 477083 23218 477125 23454
rect 476805 23134 477125 23218
rect 476805 22898 476847 23134
rect 477083 22898 477125 23134
rect 476805 22866 477125 22898
rect 498874 23454 499194 23486
rect 498874 23218 498916 23454
rect 499152 23218 499194 23454
rect 498874 23134 499194 23218
rect 498874 22898 498916 23134
rect 499152 22898 499194 23134
rect 498874 22866 499194 22898
rect 504805 23454 505125 23486
rect 504805 23218 504847 23454
rect 505083 23218 505125 23454
rect 504805 23134 505125 23218
rect 504805 22898 504847 23134
rect 505083 22898 505125 23134
rect 504805 22866 505125 22898
rect 526874 23454 527194 23486
rect 526874 23218 526916 23454
rect 527152 23218 527194 23454
rect 526874 23134 527194 23218
rect 526874 22898 526916 23134
rect 527152 22898 527194 23134
rect 526874 22866 527194 22898
rect 532805 23454 533125 23486
rect 532805 23218 532847 23454
rect 533083 23218 533125 23454
rect 532805 23134 533125 23218
rect 532805 22898 532847 23134
rect 533083 22898 533125 23134
rect 532805 22866 533125 22898
rect 554874 23454 555194 23486
rect 554874 23218 554916 23454
rect 555152 23218 555194 23454
rect 554874 23134 555194 23218
rect 554874 22898 554916 23134
rect 555152 22898 555194 23134
rect 554874 22866 555194 22898
rect 560805 23454 561125 23486
rect 560805 23218 560847 23454
rect 561083 23218 561125 23454
rect 560805 23134 561125 23218
rect 560805 22898 560847 23134
rect 561083 22898 561125 23134
rect 560805 22866 561125 22898
rect 65994 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 66614 -1306
rect 65994 -1626 66614 -1542
rect 65994 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 66614 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 65994 -7654 66614 -1862
rect 573494 -346 574114 26273
rect 573494 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 574114 -346
rect 573494 -666 574114 -582
rect 573494 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 574114 -666
rect 573494 -7654 574114 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 701829 585930 704282
rect 585310 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 585930 701829
rect 585310 701509 585930 701593
rect 585310 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 585930 701509
rect 585310 674829 585930 701273
rect 585310 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 585930 674829
rect 585310 674509 585930 674593
rect 585310 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 585930 674509
rect 585310 647829 585930 674273
rect 585310 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 585930 647829
rect 585310 647509 585930 647593
rect 585310 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 585930 647509
rect 585310 620829 585930 647273
rect 585310 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 585930 620829
rect 585310 620509 585930 620593
rect 585310 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 585930 620509
rect 585310 593829 585930 620273
rect 585310 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 585930 593829
rect 585310 593509 585930 593593
rect 585310 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 585930 593509
rect 585310 566829 585930 593273
rect 585310 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 585930 566829
rect 585310 566509 585930 566593
rect 585310 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 585930 566509
rect 585310 539829 585930 566273
rect 585310 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 585930 539829
rect 585310 539509 585930 539593
rect 585310 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 585930 539509
rect 585310 512829 585930 539273
rect 585310 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 585930 512829
rect 585310 512509 585930 512593
rect 585310 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 585930 512509
rect 585310 485829 585930 512273
rect 585310 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 585930 485829
rect 585310 485509 585930 485593
rect 585310 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 585930 485509
rect 585310 458829 585930 485273
rect 585310 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 585930 458829
rect 585310 458509 585930 458593
rect 585310 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 585930 458509
rect 585310 431829 585930 458273
rect 585310 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 585930 431829
rect 585310 431509 585930 431593
rect 585310 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 585930 431509
rect 585310 404829 585930 431273
rect 585310 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 585930 404829
rect 585310 404509 585930 404593
rect 585310 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 585930 404509
rect 585310 377829 585930 404273
rect 585310 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 585930 377829
rect 585310 377509 585930 377593
rect 585310 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 585930 377509
rect 585310 350829 585930 377273
rect 585310 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 585930 350829
rect 585310 350509 585930 350593
rect 585310 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 585930 350509
rect 585310 323829 585930 350273
rect 585310 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 585930 323829
rect 585310 323509 585930 323593
rect 585310 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 585930 323509
rect 585310 296829 585930 323273
rect 585310 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 585930 296829
rect 585310 296509 585930 296593
rect 585310 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 585930 296509
rect 585310 269829 585930 296273
rect 585310 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 585930 269829
rect 585310 269509 585930 269593
rect 585310 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 585930 269509
rect 585310 242829 585930 269273
rect 585310 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 585930 242829
rect 585310 242509 585930 242593
rect 585310 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 585930 242509
rect 585310 215829 585930 242273
rect 585310 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 585930 215829
rect 585310 215509 585930 215593
rect 585310 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 585930 215509
rect 585310 188829 585930 215273
rect 585310 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 585930 188829
rect 585310 188509 585930 188593
rect 585310 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 585930 188509
rect 585310 161829 585930 188273
rect 585310 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 585930 161829
rect 585310 161509 585930 161593
rect 585310 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 585930 161509
rect 585310 134829 585930 161273
rect 585310 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 585930 134829
rect 585310 134509 585930 134593
rect 585310 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 585930 134509
rect 585310 107829 585930 134273
rect 585310 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 585930 107829
rect 585310 107509 585930 107593
rect 585310 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 585930 107509
rect 585310 80829 585930 107273
rect 585310 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 585930 80829
rect 585310 80509 585930 80593
rect 585310 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 585930 80509
rect 585310 53829 585930 80273
rect 585310 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 585930 53829
rect 585310 53509 585930 53593
rect 585310 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 585930 53509
rect 585310 26829 585930 53273
rect 585310 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 585930 26829
rect 585310 26509 585930 26593
rect 585310 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 585930 26509
rect 585310 -346 585930 26273
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 698454 586890 705242
rect 586270 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 586890 698454
rect 586270 698134 586890 698218
rect 586270 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 586890 698134
rect 586270 671454 586890 697898
rect 586270 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 586890 671454
rect 586270 671134 586890 671218
rect 586270 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 586890 671134
rect 586270 644454 586890 670898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 617454 586890 643898
rect 586270 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 586890 617454
rect 586270 617134 586890 617218
rect 586270 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 586890 617134
rect 586270 590454 586890 616898
rect 586270 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 586890 590454
rect 586270 590134 586890 590218
rect 586270 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 586890 590134
rect 586270 563454 586890 589898
rect 586270 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 586890 563454
rect 586270 563134 586890 563218
rect 586270 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 586890 563134
rect 586270 536454 586890 562898
rect 586270 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 586890 536454
rect 586270 536134 586890 536218
rect 586270 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 586890 536134
rect 586270 509454 586890 535898
rect 586270 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 586890 509454
rect 586270 509134 586890 509218
rect 586270 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 586890 509134
rect 586270 482454 586890 508898
rect 586270 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 586890 482454
rect 586270 482134 586890 482218
rect 586270 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 586890 482134
rect 586270 455454 586890 481898
rect 586270 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 586890 455454
rect 586270 455134 586890 455218
rect 586270 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 586890 455134
rect 586270 428454 586890 454898
rect 586270 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 586890 428454
rect 586270 428134 586890 428218
rect 586270 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 586890 428134
rect 586270 401454 586890 427898
rect 586270 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 586890 401454
rect 586270 401134 586890 401218
rect 586270 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 586890 401134
rect 586270 374454 586890 400898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 347454 586890 373898
rect 586270 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 586890 347454
rect 586270 347134 586890 347218
rect 586270 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 586890 347134
rect 586270 320454 586890 346898
rect 586270 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 586890 320454
rect 586270 320134 586890 320218
rect 586270 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 586890 320134
rect 586270 293454 586890 319898
rect 586270 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 586890 293454
rect 586270 293134 586890 293218
rect 586270 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 586890 293134
rect 586270 266454 586890 292898
rect 586270 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 586890 266454
rect 586270 266134 586890 266218
rect 586270 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 586890 266134
rect 586270 239454 586890 265898
rect 586270 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 586890 239454
rect 586270 239134 586890 239218
rect 586270 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 586890 239134
rect 586270 212454 586890 238898
rect 586270 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect 586270 212134 586890 212218
rect 586270 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect 586270 185454 586890 211898
rect 586270 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 586890 185454
rect 586270 185134 586890 185218
rect 586270 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 586890 185134
rect 586270 158454 586890 184898
rect 586270 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 586890 158454
rect 586270 158134 586890 158218
rect 586270 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 586890 158134
rect 586270 131454 586890 157898
rect 586270 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 586890 131454
rect 586270 131134 586890 131218
rect 586270 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 586890 131134
rect 586270 104454 586890 130898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 77454 586890 103898
rect 586270 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 586890 77454
rect 586270 77134 586890 77218
rect 586270 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 586890 77134
rect 586270 50454 586890 76898
rect 586270 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 586890 50454
rect 586270 50134 586890 50218
rect 586270 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 586890 50134
rect 586270 23454 586890 49898
rect 586270 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 586890 23454
rect 586270 23134 586890 23218
rect 586270 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 586890 23134
rect 586270 -1306 586890 22898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 38026 705562 38262 705798
rect 38346 705562 38582 705798
rect 38026 705242 38262 705478
rect 38346 705242 38582 705478
rect -2934 698218 -2698 698454
rect -2614 698218 -2378 698454
rect -2934 697898 -2698 698134
rect -2614 697898 -2378 698134
rect -2934 671218 -2698 671454
rect -2614 671218 -2378 671454
rect -2934 670898 -2698 671134
rect -2614 670898 -2378 671134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 617218 -2698 617454
rect -2614 617218 -2378 617454
rect -2934 616898 -2698 617134
rect -2614 616898 -2378 617134
rect -2934 590218 -2698 590454
rect -2614 590218 -2378 590454
rect -2934 589898 -2698 590134
rect -2614 589898 -2378 590134
rect -2934 563218 -2698 563454
rect -2614 563218 -2378 563454
rect -2934 562898 -2698 563134
rect -2614 562898 -2378 563134
rect -2934 536218 -2698 536454
rect -2614 536218 -2378 536454
rect -2934 535898 -2698 536134
rect -2614 535898 -2378 536134
rect -2934 509218 -2698 509454
rect -2614 509218 -2378 509454
rect -2934 508898 -2698 509134
rect -2614 508898 -2378 509134
rect -2934 482218 -2698 482454
rect -2614 482218 -2378 482454
rect -2934 481898 -2698 482134
rect -2614 481898 -2378 482134
rect -2934 455218 -2698 455454
rect -2614 455218 -2378 455454
rect -2934 454898 -2698 455134
rect -2614 454898 -2378 455134
rect -2934 428218 -2698 428454
rect -2614 428218 -2378 428454
rect -2934 427898 -2698 428134
rect -2614 427898 -2378 428134
rect -2934 401218 -2698 401454
rect -2614 401218 -2378 401454
rect -2934 400898 -2698 401134
rect -2614 400898 -2378 401134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 347218 -2698 347454
rect -2614 347218 -2378 347454
rect -2934 346898 -2698 347134
rect -2614 346898 -2378 347134
rect -2934 320218 -2698 320454
rect -2614 320218 -2378 320454
rect -2934 319898 -2698 320134
rect -2614 319898 -2378 320134
rect -2934 293218 -2698 293454
rect -2614 293218 -2378 293454
rect -2934 292898 -2698 293134
rect -2614 292898 -2378 293134
rect -2934 266218 -2698 266454
rect -2614 266218 -2378 266454
rect -2934 265898 -2698 266134
rect -2614 265898 -2378 266134
rect -2934 239218 -2698 239454
rect -2614 239218 -2378 239454
rect -2934 238898 -2698 239134
rect -2614 238898 -2378 239134
rect -2934 212218 -2698 212454
rect -2614 212218 -2378 212454
rect -2934 211898 -2698 212134
rect -2614 211898 -2378 212134
rect -2934 185218 -2698 185454
rect -2614 185218 -2378 185454
rect -2934 184898 -2698 185134
rect -2614 184898 -2378 185134
rect -2934 158218 -2698 158454
rect -2614 158218 -2378 158454
rect -2934 157898 -2698 158134
rect -2614 157898 -2378 158134
rect -2934 131218 -2698 131454
rect -2614 131218 -2378 131454
rect -2934 130898 -2698 131134
rect -2614 130898 -2378 131134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 77218 -2698 77454
rect -2614 77218 -2378 77454
rect -2934 76898 -2698 77134
rect -2614 76898 -2378 77134
rect -2934 50218 -2698 50454
rect -2614 50218 -2378 50454
rect -2934 49898 -2698 50134
rect -2614 49898 -2378 50134
rect -2934 23218 -2698 23454
rect -2614 23218 -2378 23454
rect -2934 22898 -2698 23134
rect -2614 22898 -2378 23134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 701593 -1738 701829
rect -1654 701593 -1418 701829
rect -1974 701273 -1738 701509
rect -1654 701273 -1418 701509
rect 38026 698218 38262 698454
rect 38346 698218 38582 698454
rect 38026 697898 38262 698134
rect 38346 697898 38582 698134
rect 41526 704602 41762 704838
rect 41846 704602 42082 704838
rect 41526 704282 41762 704518
rect 41846 704282 42082 704518
rect 41526 701593 41762 701829
rect 41846 701593 42082 701829
rect 41526 701273 41762 701509
rect 41846 701273 42082 701509
rect 66026 705562 66262 705798
rect 66346 705562 66582 705798
rect 66026 705242 66262 705478
rect 66346 705242 66582 705478
rect 66026 698218 66262 698454
rect 66346 698218 66582 698454
rect 66026 697898 66262 698134
rect 66346 697898 66582 698134
rect 69526 704602 69762 704838
rect 69846 704602 70082 704838
rect 69526 704282 69762 704518
rect 69846 704282 70082 704518
rect 69526 701593 69762 701829
rect 69846 701593 70082 701829
rect 69526 701273 69762 701509
rect 69846 701273 70082 701509
rect 94026 705562 94262 705798
rect 94346 705562 94582 705798
rect 94026 705242 94262 705478
rect 94346 705242 94582 705478
rect 94026 698218 94262 698454
rect 94346 698218 94582 698454
rect 94026 697898 94262 698134
rect 94346 697898 94582 698134
rect 97526 704602 97762 704838
rect 97846 704602 98082 704838
rect 97526 704282 97762 704518
rect 97846 704282 98082 704518
rect 97526 701593 97762 701829
rect 97846 701593 98082 701829
rect 97526 701273 97762 701509
rect 97846 701273 98082 701509
rect 122026 705562 122262 705798
rect 122346 705562 122582 705798
rect 122026 705242 122262 705478
rect 122346 705242 122582 705478
rect 122026 698218 122262 698454
rect 122346 698218 122582 698454
rect 122026 697898 122262 698134
rect 122346 697898 122582 698134
rect 125526 704602 125762 704838
rect 125846 704602 126082 704838
rect 125526 704282 125762 704518
rect 125846 704282 126082 704518
rect 125526 701593 125762 701829
rect 125846 701593 126082 701829
rect 125526 701273 125762 701509
rect 125846 701273 126082 701509
rect 150026 705562 150262 705798
rect 150346 705562 150582 705798
rect 150026 705242 150262 705478
rect 150346 705242 150582 705478
rect 150026 698218 150262 698454
rect 150346 698218 150582 698454
rect 150026 697898 150262 698134
rect 150346 697898 150582 698134
rect 153526 704602 153762 704838
rect 153846 704602 154082 704838
rect 153526 704282 153762 704518
rect 153846 704282 154082 704518
rect 153526 701593 153762 701829
rect 153846 701593 154082 701829
rect 153526 701273 153762 701509
rect 153846 701273 154082 701509
rect 178026 705562 178262 705798
rect 178346 705562 178582 705798
rect 178026 705242 178262 705478
rect 178346 705242 178582 705478
rect 178026 698218 178262 698454
rect 178346 698218 178582 698454
rect 178026 697898 178262 698134
rect 178346 697898 178582 698134
rect 181526 704602 181762 704838
rect 181846 704602 182082 704838
rect 181526 704282 181762 704518
rect 181846 704282 182082 704518
rect 181526 701593 181762 701829
rect 181846 701593 182082 701829
rect 181526 701273 181762 701509
rect 181846 701273 182082 701509
rect 206026 705562 206262 705798
rect 206346 705562 206582 705798
rect 206026 705242 206262 705478
rect 206346 705242 206582 705478
rect 206026 698218 206262 698454
rect 206346 698218 206582 698454
rect 206026 697898 206262 698134
rect 206346 697898 206582 698134
rect 209526 704602 209762 704838
rect 209846 704602 210082 704838
rect 209526 704282 209762 704518
rect 209846 704282 210082 704518
rect 209526 701593 209762 701829
rect 209846 701593 210082 701829
rect 209526 701273 209762 701509
rect 209846 701273 210082 701509
rect 234026 705562 234262 705798
rect 234346 705562 234582 705798
rect 234026 705242 234262 705478
rect 234346 705242 234582 705478
rect 234026 698218 234262 698454
rect 234346 698218 234582 698454
rect 234026 697898 234262 698134
rect 234346 697898 234582 698134
rect 237526 704602 237762 704838
rect 237846 704602 238082 704838
rect 237526 704282 237762 704518
rect 237846 704282 238082 704518
rect 237526 701593 237762 701829
rect 237846 701593 238082 701829
rect 237526 701273 237762 701509
rect 237846 701273 238082 701509
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 262026 698218 262262 698454
rect 262346 698218 262582 698454
rect 262026 697898 262262 698134
rect 262346 697898 262582 698134
rect 265526 704602 265762 704838
rect 265846 704602 266082 704838
rect 265526 704282 265762 704518
rect 265846 704282 266082 704518
rect 265526 701593 265762 701829
rect 265846 701593 266082 701829
rect 265526 701273 265762 701509
rect 265846 701273 266082 701509
rect 290026 705562 290262 705798
rect 290346 705562 290582 705798
rect 290026 705242 290262 705478
rect 290346 705242 290582 705478
rect 290026 698218 290262 698454
rect 290346 698218 290582 698454
rect 290026 697898 290262 698134
rect 290346 697898 290582 698134
rect 293526 704602 293762 704838
rect 293846 704602 294082 704838
rect 293526 704282 293762 704518
rect 293846 704282 294082 704518
rect 293526 701593 293762 701829
rect 293846 701593 294082 701829
rect 293526 701273 293762 701509
rect 293846 701273 294082 701509
rect 318026 705562 318262 705798
rect 318346 705562 318582 705798
rect 318026 705242 318262 705478
rect 318346 705242 318582 705478
rect 318026 698218 318262 698454
rect 318346 698218 318582 698454
rect 318026 697898 318262 698134
rect 318346 697898 318582 698134
rect 321526 704602 321762 704838
rect 321846 704602 322082 704838
rect 321526 704282 321762 704518
rect 321846 704282 322082 704518
rect 321526 701593 321762 701829
rect 321846 701593 322082 701829
rect 321526 701273 321762 701509
rect 321846 701273 322082 701509
rect 346026 705562 346262 705798
rect 346346 705562 346582 705798
rect 346026 705242 346262 705478
rect 346346 705242 346582 705478
rect 346026 698218 346262 698454
rect 346346 698218 346582 698454
rect 346026 697898 346262 698134
rect 346346 697898 346582 698134
rect 349526 704602 349762 704838
rect 349846 704602 350082 704838
rect 349526 704282 349762 704518
rect 349846 704282 350082 704518
rect 349526 701593 349762 701829
rect 349846 701593 350082 701829
rect 349526 701273 349762 701509
rect 349846 701273 350082 701509
rect 374026 705562 374262 705798
rect 374346 705562 374582 705798
rect 374026 705242 374262 705478
rect 374346 705242 374582 705478
rect 374026 698218 374262 698454
rect 374346 698218 374582 698454
rect 374026 697898 374262 698134
rect 374346 697898 374582 698134
rect 377526 704602 377762 704838
rect 377846 704602 378082 704838
rect 377526 704282 377762 704518
rect 377846 704282 378082 704518
rect 377526 701593 377762 701829
rect 377846 701593 378082 701829
rect 377526 701273 377762 701509
rect 377846 701273 378082 701509
rect 402026 705562 402262 705798
rect 402346 705562 402582 705798
rect 402026 705242 402262 705478
rect 402346 705242 402582 705478
rect 402026 698218 402262 698454
rect 402346 698218 402582 698454
rect 402026 697898 402262 698134
rect 402346 697898 402582 698134
rect 405526 704602 405762 704838
rect 405846 704602 406082 704838
rect 405526 704282 405762 704518
rect 405846 704282 406082 704518
rect 405526 701593 405762 701829
rect 405846 701593 406082 701829
rect 405526 701273 405762 701509
rect 405846 701273 406082 701509
rect 430026 705562 430262 705798
rect 430346 705562 430582 705798
rect 430026 705242 430262 705478
rect 430346 705242 430582 705478
rect 430026 698218 430262 698454
rect 430346 698218 430582 698454
rect 430026 697898 430262 698134
rect 430346 697898 430582 698134
rect 433526 704602 433762 704838
rect 433846 704602 434082 704838
rect 433526 704282 433762 704518
rect 433846 704282 434082 704518
rect 433526 701593 433762 701829
rect 433846 701593 434082 701829
rect 433526 701273 433762 701509
rect 433846 701273 434082 701509
rect 458026 705562 458262 705798
rect 458346 705562 458582 705798
rect 458026 705242 458262 705478
rect 458346 705242 458582 705478
rect 458026 698218 458262 698454
rect 458346 698218 458582 698454
rect 458026 697898 458262 698134
rect 458346 697898 458582 698134
rect 461526 704602 461762 704838
rect 461846 704602 462082 704838
rect 461526 704282 461762 704518
rect 461846 704282 462082 704518
rect 461526 701593 461762 701829
rect 461846 701593 462082 701829
rect 461526 701273 461762 701509
rect 461846 701273 462082 701509
rect 486026 705562 486262 705798
rect 486346 705562 486582 705798
rect 486026 705242 486262 705478
rect 486346 705242 486582 705478
rect 486026 698218 486262 698454
rect 486346 698218 486582 698454
rect 486026 697898 486262 698134
rect 486346 697898 486582 698134
rect 489526 704602 489762 704838
rect 489846 704602 490082 704838
rect 489526 704282 489762 704518
rect 489846 704282 490082 704518
rect 489526 701593 489762 701829
rect 489846 701593 490082 701829
rect 489526 701273 489762 701509
rect 489846 701273 490082 701509
rect 514026 705562 514262 705798
rect 514346 705562 514582 705798
rect 514026 705242 514262 705478
rect 514346 705242 514582 705478
rect 514026 698218 514262 698454
rect 514346 698218 514582 698454
rect 514026 697898 514262 698134
rect 514346 697898 514582 698134
rect 517526 704602 517762 704838
rect 517846 704602 518082 704838
rect 517526 704282 517762 704518
rect 517846 704282 518082 704518
rect 517526 701593 517762 701829
rect 517846 701593 518082 701829
rect 517526 701273 517762 701509
rect 517846 701273 518082 701509
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 542026 698218 542262 698454
rect 542346 698218 542582 698454
rect 542026 697898 542262 698134
rect 542346 697898 542582 698134
rect 545526 704602 545762 704838
rect 545846 704602 546082 704838
rect 545526 704282 545762 704518
rect 545846 704282 546082 704518
rect 545526 701593 545762 701829
rect 545846 701593 546082 701829
rect 545526 701273 545762 701509
rect 545846 701273 546082 701509
rect 570026 705562 570262 705798
rect 570346 705562 570582 705798
rect 570026 705242 570262 705478
rect 570346 705242 570582 705478
rect 570026 698218 570262 698454
rect 570346 698218 570582 698454
rect 570026 697898 570262 698134
rect 570346 697898 570582 698134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 573526 704602 573762 704838
rect 573846 704602 574082 704838
rect 573526 704282 573762 704518
rect 573846 704282 574082 704518
rect 573526 701593 573762 701829
rect 573846 701593 574082 701829
rect 573526 701273 573762 701509
rect 573846 701273 574082 701509
rect -1974 674593 -1738 674829
rect -1654 674593 -1418 674829
rect -1974 674273 -1738 674509
rect -1654 674273 -1418 674509
rect 19952 674593 20188 674829
rect 19952 674273 20188 674509
rect 25882 674593 26118 674829
rect 25882 674273 26118 674509
rect 31813 674593 32049 674829
rect 31813 674273 32049 674509
rect 47952 674593 48188 674829
rect 47952 674273 48188 674509
rect 53882 674593 54118 674829
rect 53882 674273 54118 674509
rect 59813 674593 60049 674829
rect 59813 674273 60049 674509
rect 75952 674593 76188 674829
rect 75952 674273 76188 674509
rect 81882 674593 82118 674829
rect 81882 674273 82118 674509
rect 87813 674593 88049 674829
rect 87813 674273 88049 674509
rect 103952 674593 104188 674829
rect 103952 674273 104188 674509
rect 109882 674593 110118 674829
rect 109882 674273 110118 674509
rect 115813 674593 116049 674829
rect 115813 674273 116049 674509
rect 131952 674593 132188 674829
rect 131952 674273 132188 674509
rect 137882 674593 138118 674829
rect 137882 674273 138118 674509
rect 143813 674593 144049 674829
rect 143813 674273 144049 674509
rect 159952 674593 160188 674829
rect 159952 674273 160188 674509
rect 165882 674593 166118 674829
rect 165882 674273 166118 674509
rect 171813 674593 172049 674829
rect 171813 674273 172049 674509
rect 187952 674593 188188 674829
rect 187952 674273 188188 674509
rect 193882 674593 194118 674829
rect 193882 674273 194118 674509
rect 199813 674593 200049 674829
rect 199813 674273 200049 674509
rect 215952 674593 216188 674829
rect 215952 674273 216188 674509
rect 221882 674593 222118 674829
rect 221882 674273 222118 674509
rect 227813 674593 228049 674829
rect 227813 674273 228049 674509
rect 243952 674593 244188 674829
rect 243952 674273 244188 674509
rect 249882 674593 250118 674829
rect 249882 674273 250118 674509
rect 255813 674593 256049 674829
rect 255813 674273 256049 674509
rect 271952 674593 272188 674829
rect 271952 674273 272188 674509
rect 277882 674593 278118 674829
rect 277882 674273 278118 674509
rect 283813 674593 284049 674829
rect 283813 674273 284049 674509
rect 299952 674593 300188 674829
rect 299952 674273 300188 674509
rect 305882 674593 306118 674829
rect 305882 674273 306118 674509
rect 311813 674593 312049 674829
rect 311813 674273 312049 674509
rect 327952 674593 328188 674829
rect 327952 674273 328188 674509
rect 333882 674593 334118 674829
rect 333882 674273 334118 674509
rect 339813 674593 340049 674829
rect 339813 674273 340049 674509
rect 355952 674593 356188 674829
rect 355952 674273 356188 674509
rect 361882 674593 362118 674829
rect 361882 674273 362118 674509
rect 367813 674593 368049 674829
rect 367813 674273 368049 674509
rect 383952 674593 384188 674829
rect 383952 674273 384188 674509
rect 389882 674593 390118 674829
rect 389882 674273 390118 674509
rect 395813 674593 396049 674829
rect 395813 674273 396049 674509
rect 411952 674593 412188 674829
rect 411952 674273 412188 674509
rect 417882 674593 418118 674829
rect 417882 674273 418118 674509
rect 423813 674593 424049 674829
rect 423813 674273 424049 674509
rect 439952 674593 440188 674829
rect 439952 674273 440188 674509
rect 445882 674593 446118 674829
rect 445882 674273 446118 674509
rect 451813 674593 452049 674829
rect 451813 674273 452049 674509
rect 467952 674593 468188 674829
rect 467952 674273 468188 674509
rect 473882 674593 474118 674829
rect 473882 674273 474118 674509
rect 479813 674593 480049 674829
rect 479813 674273 480049 674509
rect 495952 674593 496188 674829
rect 495952 674273 496188 674509
rect 501882 674593 502118 674829
rect 501882 674273 502118 674509
rect 507813 674593 508049 674829
rect 507813 674273 508049 674509
rect 523952 674593 524188 674829
rect 523952 674273 524188 674509
rect 529882 674593 530118 674829
rect 529882 674273 530118 674509
rect 535813 674593 536049 674829
rect 535813 674273 536049 674509
rect 551952 674593 552188 674829
rect 551952 674273 552188 674509
rect 557882 674593 558118 674829
rect 557882 674273 558118 674509
rect 563813 674593 564049 674829
rect 563813 674273 564049 674509
rect 573526 674593 573762 674829
rect 573846 674593 574082 674829
rect 573526 674273 573762 674509
rect 573846 674273 574082 674509
rect 22916 671218 23152 671454
rect 22916 670898 23152 671134
rect 28847 671218 29083 671454
rect 28847 670898 29083 671134
rect 50916 671218 51152 671454
rect 50916 670898 51152 671134
rect 56847 671218 57083 671454
rect 56847 670898 57083 671134
rect 78916 671218 79152 671454
rect 78916 670898 79152 671134
rect 84847 671218 85083 671454
rect 84847 670898 85083 671134
rect 106916 671218 107152 671454
rect 106916 670898 107152 671134
rect 112847 671218 113083 671454
rect 112847 670898 113083 671134
rect 134916 671218 135152 671454
rect 134916 670898 135152 671134
rect 140847 671218 141083 671454
rect 140847 670898 141083 671134
rect 162916 671218 163152 671454
rect 162916 670898 163152 671134
rect 168847 671218 169083 671454
rect 168847 670898 169083 671134
rect 190916 671218 191152 671454
rect 190916 670898 191152 671134
rect 196847 671218 197083 671454
rect 196847 670898 197083 671134
rect 218916 671218 219152 671454
rect 218916 670898 219152 671134
rect 224847 671218 225083 671454
rect 224847 670898 225083 671134
rect 246916 671218 247152 671454
rect 246916 670898 247152 671134
rect 252847 671218 253083 671454
rect 252847 670898 253083 671134
rect 274916 671218 275152 671454
rect 274916 670898 275152 671134
rect 280847 671218 281083 671454
rect 280847 670898 281083 671134
rect 302916 671218 303152 671454
rect 302916 670898 303152 671134
rect 308847 671218 309083 671454
rect 308847 670898 309083 671134
rect 330916 671218 331152 671454
rect 330916 670898 331152 671134
rect 336847 671218 337083 671454
rect 336847 670898 337083 671134
rect 358916 671218 359152 671454
rect 358916 670898 359152 671134
rect 364847 671218 365083 671454
rect 364847 670898 365083 671134
rect 386916 671218 387152 671454
rect 386916 670898 387152 671134
rect 392847 671218 393083 671454
rect 392847 670898 393083 671134
rect 414916 671218 415152 671454
rect 414916 670898 415152 671134
rect 420847 671218 421083 671454
rect 420847 670898 421083 671134
rect 442916 671218 443152 671454
rect 442916 670898 443152 671134
rect 448847 671218 449083 671454
rect 448847 670898 449083 671134
rect 470916 671218 471152 671454
rect 470916 670898 471152 671134
rect 476847 671218 477083 671454
rect 476847 670898 477083 671134
rect 498916 671218 499152 671454
rect 498916 670898 499152 671134
rect 504847 671218 505083 671454
rect 504847 670898 505083 671134
rect 526916 671218 527152 671454
rect 526916 670898 527152 671134
rect 532847 671218 533083 671454
rect 532847 670898 533083 671134
rect 554916 671218 555152 671454
rect 554916 670898 555152 671134
rect 560847 671218 561083 671454
rect 560847 670898 561083 671134
rect -1974 647593 -1738 647829
rect -1654 647593 -1418 647829
rect -1974 647273 -1738 647509
rect -1654 647273 -1418 647509
rect 19952 647593 20188 647829
rect 19952 647273 20188 647509
rect 25882 647593 26118 647829
rect 25882 647273 26118 647509
rect 31813 647593 32049 647829
rect 31813 647273 32049 647509
rect 47952 647593 48188 647829
rect 47952 647273 48188 647509
rect 53882 647593 54118 647829
rect 53882 647273 54118 647509
rect 59813 647593 60049 647829
rect 59813 647273 60049 647509
rect 75952 647593 76188 647829
rect 75952 647273 76188 647509
rect 81882 647593 82118 647829
rect 81882 647273 82118 647509
rect 87813 647593 88049 647829
rect 87813 647273 88049 647509
rect 103952 647593 104188 647829
rect 103952 647273 104188 647509
rect 109882 647593 110118 647829
rect 109882 647273 110118 647509
rect 115813 647593 116049 647829
rect 115813 647273 116049 647509
rect 131952 647593 132188 647829
rect 131952 647273 132188 647509
rect 137882 647593 138118 647829
rect 137882 647273 138118 647509
rect 143813 647593 144049 647829
rect 143813 647273 144049 647509
rect 159952 647593 160188 647829
rect 159952 647273 160188 647509
rect 165882 647593 166118 647829
rect 165882 647273 166118 647509
rect 171813 647593 172049 647829
rect 171813 647273 172049 647509
rect 187952 647593 188188 647829
rect 187952 647273 188188 647509
rect 193882 647593 194118 647829
rect 193882 647273 194118 647509
rect 199813 647593 200049 647829
rect 199813 647273 200049 647509
rect 215952 647593 216188 647829
rect 215952 647273 216188 647509
rect 221882 647593 222118 647829
rect 221882 647273 222118 647509
rect 227813 647593 228049 647829
rect 227813 647273 228049 647509
rect 243952 647593 244188 647829
rect 243952 647273 244188 647509
rect 249882 647593 250118 647829
rect 249882 647273 250118 647509
rect 255813 647593 256049 647829
rect 255813 647273 256049 647509
rect 271952 647593 272188 647829
rect 271952 647273 272188 647509
rect 277882 647593 278118 647829
rect 277882 647273 278118 647509
rect 283813 647593 284049 647829
rect 283813 647273 284049 647509
rect 299952 647593 300188 647829
rect 299952 647273 300188 647509
rect 305882 647593 306118 647829
rect 305882 647273 306118 647509
rect 311813 647593 312049 647829
rect 311813 647273 312049 647509
rect 327952 647593 328188 647829
rect 327952 647273 328188 647509
rect 333882 647593 334118 647829
rect 333882 647273 334118 647509
rect 339813 647593 340049 647829
rect 339813 647273 340049 647509
rect 355952 647593 356188 647829
rect 355952 647273 356188 647509
rect 361882 647593 362118 647829
rect 361882 647273 362118 647509
rect 367813 647593 368049 647829
rect 367813 647273 368049 647509
rect 383952 647593 384188 647829
rect 383952 647273 384188 647509
rect 389882 647593 390118 647829
rect 389882 647273 390118 647509
rect 395813 647593 396049 647829
rect 395813 647273 396049 647509
rect 411952 647593 412188 647829
rect 411952 647273 412188 647509
rect 417882 647593 418118 647829
rect 417882 647273 418118 647509
rect 423813 647593 424049 647829
rect 423813 647273 424049 647509
rect 439952 647593 440188 647829
rect 439952 647273 440188 647509
rect 445882 647593 446118 647829
rect 445882 647273 446118 647509
rect 451813 647593 452049 647829
rect 451813 647273 452049 647509
rect 467952 647593 468188 647829
rect 467952 647273 468188 647509
rect 473882 647593 474118 647829
rect 473882 647273 474118 647509
rect 479813 647593 480049 647829
rect 479813 647273 480049 647509
rect 495952 647593 496188 647829
rect 495952 647273 496188 647509
rect 501882 647593 502118 647829
rect 501882 647273 502118 647509
rect 507813 647593 508049 647829
rect 507813 647273 508049 647509
rect 523952 647593 524188 647829
rect 523952 647273 524188 647509
rect 529882 647593 530118 647829
rect 529882 647273 530118 647509
rect 535813 647593 536049 647829
rect 535813 647273 536049 647509
rect 551952 647593 552188 647829
rect 551952 647273 552188 647509
rect 557882 647593 558118 647829
rect 557882 647273 558118 647509
rect 563813 647593 564049 647829
rect 563813 647273 564049 647509
rect 573526 647593 573762 647829
rect 573846 647593 574082 647829
rect 573526 647273 573762 647509
rect 573846 647273 574082 647509
rect 22916 644218 23152 644454
rect 22916 643898 23152 644134
rect 28847 644218 29083 644454
rect 28847 643898 29083 644134
rect 50916 644218 51152 644454
rect 50916 643898 51152 644134
rect 56847 644218 57083 644454
rect 56847 643898 57083 644134
rect 78916 644218 79152 644454
rect 78916 643898 79152 644134
rect 84847 644218 85083 644454
rect 84847 643898 85083 644134
rect 106916 644218 107152 644454
rect 106916 643898 107152 644134
rect 112847 644218 113083 644454
rect 112847 643898 113083 644134
rect 134916 644218 135152 644454
rect 134916 643898 135152 644134
rect 140847 644218 141083 644454
rect 140847 643898 141083 644134
rect 162916 644218 163152 644454
rect 162916 643898 163152 644134
rect 168847 644218 169083 644454
rect 168847 643898 169083 644134
rect 190916 644218 191152 644454
rect 190916 643898 191152 644134
rect 196847 644218 197083 644454
rect 196847 643898 197083 644134
rect 218916 644218 219152 644454
rect 218916 643898 219152 644134
rect 224847 644218 225083 644454
rect 224847 643898 225083 644134
rect 246916 644218 247152 644454
rect 246916 643898 247152 644134
rect 252847 644218 253083 644454
rect 252847 643898 253083 644134
rect 274916 644218 275152 644454
rect 274916 643898 275152 644134
rect 280847 644218 281083 644454
rect 280847 643898 281083 644134
rect 302916 644218 303152 644454
rect 302916 643898 303152 644134
rect 308847 644218 309083 644454
rect 308847 643898 309083 644134
rect 330916 644218 331152 644454
rect 330916 643898 331152 644134
rect 336847 644218 337083 644454
rect 336847 643898 337083 644134
rect 358916 644218 359152 644454
rect 358916 643898 359152 644134
rect 364847 644218 365083 644454
rect 364847 643898 365083 644134
rect 386916 644218 387152 644454
rect 386916 643898 387152 644134
rect 392847 644218 393083 644454
rect 392847 643898 393083 644134
rect 414916 644218 415152 644454
rect 414916 643898 415152 644134
rect 420847 644218 421083 644454
rect 420847 643898 421083 644134
rect 442916 644218 443152 644454
rect 442916 643898 443152 644134
rect 448847 644218 449083 644454
rect 448847 643898 449083 644134
rect 470916 644218 471152 644454
rect 470916 643898 471152 644134
rect 476847 644218 477083 644454
rect 476847 643898 477083 644134
rect 498916 644218 499152 644454
rect 498916 643898 499152 644134
rect 504847 644218 505083 644454
rect 504847 643898 505083 644134
rect 526916 644218 527152 644454
rect 526916 643898 527152 644134
rect 532847 644218 533083 644454
rect 532847 643898 533083 644134
rect 554916 644218 555152 644454
rect 554916 643898 555152 644134
rect 560847 644218 561083 644454
rect 560847 643898 561083 644134
rect -1974 620593 -1738 620829
rect -1654 620593 -1418 620829
rect -1974 620273 -1738 620509
rect -1654 620273 -1418 620509
rect 19952 620593 20188 620829
rect 19952 620273 20188 620509
rect 25882 620593 26118 620829
rect 25882 620273 26118 620509
rect 31813 620593 32049 620829
rect 31813 620273 32049 620509
rect 47952 620593 48188 620829
rect 47952 620273 48188 620509
rect 53882 620593 54118 620829
rect 53882 620273 54118 620509
rect 59813 620593 60049 620829
rect 59813 620273 60049 620509
rect 75952 620593 76188 620829
rect 75952 620273 76188 620509
rect 81882 620593 82118 620829
rect 81882 620273 82118 620509
rect 87813 620593 88049 620829
rect 87813 620273 88049 620509
rect 103952 620593 104188 620829
rect 103952 620273 104188 620509
rect 109882 620593 110118 620829
rect 109882 620273 110118 620509
rect 115813 620593 116049 620829
rect 115813 620273 116049 620509
rect 131952 620593 132188 620829
rect 131952 620273 132188 620509
rect 137882 620593 138118 620829
rect 137882 620273 138118 620509
rect 143813 620593 144049 620829
rect 143813 620273 144049 620509
rect 159952 620593 160188 620829
rect 159952 620273 160188 620509
rect 165882 620593 166118 620829
rect 165882 620273 166118 620509
rect 171813 620593 172049 620829
rect 171813 620273 172049 620509
rect 187952 620593 188188 620829
rect 187952 620273 188188 620509
rect 193882 620593 194118 620829
rect 193882 620273 194118 620509
rect 199813 620593 200049 620829
rect 199813 620273 200049 620509
rect 215952 620593 216188 620829
rect 215952 620273 216188 620509
rect 221882 620593 222118 620829
rect 221882 620273 222118 620509
rect 227813 620593 228049 620829
rect 227813 620273 228049 620509
rect 243952 620593 244188 620829
rect 243952 620273 244188 620509
rect 249882 620593 250118 620829
rect 249882 620273 250118 620509
rect 255813 620593 256049 620829
rect 255813 620273 256049 620509
rect 271952 620593 272188 620829
rect 271952 620273 272188 620509
rect 277882 620593 278118 620829
rect 277882 620273 278118 620509
rect 283813 620593 284049 620829
rect 283813 620273 284049 620509
rect 299952 620593 300188 620829
rect 299952 620273 300188 620509
rect 305882 620593 306118 620829
rect 305882 620273 306118 620509
rect 311813 620593 312049 620829
rect 311813 620273 312049 620509
rect 327952 620593 328188 620829
rect 327952 620273 328188 620509
rect 333882 620593 334118 620829
rect 333882 620273 334118 620509
rect 339813 620593 340049 620829
rect 339813 620273 340049 620509
rect 355952 620593 356188 620829
rect 355952 620273 356188 620509
rect 361882 620593 362118 620829
rect 361882 620273 362118 620509
rect 367813 620593 368049 620829
rect 367813 620273 368049 620509
rect 383952 620593 384188 620829
rect 383952 620273 384188 620509
rect 389882 620593 390118 620829
rect 389882 620273 390118 620509
rect 395813 620593 396049 620829
rect 395813 620273 396049 620509
rect 411952 620593 412188 620829
rect 411952 620273 412188 620509
rect 417882 620593 418118 620829
rect 417882 620273 418118 620509
rect 423813 620593 424049 620829
rect 423813 620273 424049 620509
rect 439952 620593 440188 620829
rect 439952 620273 440188 620509
rect 445882 620593 446118 620829
rect 445882 620273 446118 620509
rect 451813 620593 452049 620829
rect 451813 620273 452049 620509
rect 467952 620593 468188 620829
rect 467952 620273 468188 620509
rect 473882 620593 474118 620829
rect 473882 620273 474118 620509
rect 479813 620593 480049 620829
rect 479813 620273 480049 620509
rect 495952 620593 496188 620829
rect 495952 620273 496188 620509
rect 501882 620593 502118 620829
rect 501882 620273 502118 620509
rect 507813 620593 508049 620829
rect 507813 620273 508049 620509
rect 523952 620593 524188 620829
rect 523952 620273 524188 620509
rect 529882 620593 530118 620829
rect 529882 620273 530118 620509
rect 535813 620593 536049 620829
rect 535813 620273 536049 620509
rect 551952 620593 552188 620829
rect 551952 620273 552188 620509
rect 557882 620593 558118 620829
rect 557882 620273 558118 620509
rect 563813 620593 564049 620829
rect 563813 620273 564049 620509
rect 573526 620593 573762 620829
rect 573846 620593 574082 620829
rect 573526 620273 573762 620509
rect 573846 620273 574082 620509
rect 22916 617218 23152 617454
rect 22916 616898 23152 617134
rect 28847 617218 29083 617454
rect 28847 616898 29083 617134
rect 50916 617218 51152 617454
rect 50916 616898 51152 617134
rect 56847 617218 57083 617454
rect 56847 616898 57083 617134
rect 78916 617218 79152 617454
rect 78916 616898 79152 617134
rect 84847 617218 85083 617454
rect 84847 616898 85083 617134
rect 106916 617218 107152 617454
rect 106916 616898 107152 617134
rect 112847 617218 113083 617454
rect 112847 616898 113083 617134
rect 134916 617218 135152 617454
rect 134916 616898 135152 617134
rect 140847 617218 141083 617454
rect 140847 616898 141083 617134
rect 162916 617218 163152 617454
rect 162916 616898 163152 617134
rect 168847 617218 169083 617454
rect 168847 616898 169083 617134
rect 190916 617218 191152 617454
rect 190916 616898 191152 617134
rect 196847 617218 197083 617454
rect 196847 616898 197083 617134
rect 218916 617218 219152 617454
rect 218916 616898 219152 617134
rect 224847 617218 225083 617454
rect 224847 616898 225083 617134
rect 246916 617218 247152 617454
rect 246916 616898 247152 617134
rect 252847 617218 253083 617454
rect 252847 616898 253083 617134
rect 274916 617218 275152 617454
rect 274916 616898 275152 617134
rect 280847 617218 281083 617454
rect 280847 616898 281083 617134
rect 302916 617218 303152 617454
rect 302916 616898 303152 617134
rect 308847 617218 309083 617454
rect 308847 616898 309083 617134
rect 330916 617218 331152 617454
rect 330916 616898 331152 617134
rect 336847 617218 337083 617454
rect 336847 616898 337083 617134
rect 358916 617218 359152 617454
rect 358916 616898 359152 617134
rect 364847 617218 365083 617454
rect 364847 616898 365083 617134
rect 386916 617218 387152 617454
rect 386916 616898 387152 617134
rect 392847 617218 393083 617454
rect 392847 616898 393083 617134
rect 414916 617218 415152 617454
rect 414916 616898 415152 617134
rect 420847 617218 421083 617454
rect 420847 616898 421083 617134
rect 442916 617218 443152 617454
rect 442916 616898 443152 617134
rect 448847 617218 449083 617454
rect 448847 616898 449083 617134
rect 470916 617218 471152 617454
rect 470916 616898 471152 617134
rect 476847 617218 477083 617454
rect 476847 616898 477083 617134
rect 498916 617218 499152 617454
rect 498916 616898 499152 617134
rect 504847 617218 505083 617454
rect 504847 616898 505083 617134
rect 526916 617218 527152 617454
rect 526916 616898 527152 617134
rect 532847 617218 533083 617454
rect 532847 616898 533083 617134
rect 554916 617218 555152 617454
rect 554916 616898 555152 617134
rect 560847 617218 561083 617454
rect 560847 616898 561083 617134
rect -1974 593593 -1738 593829
rect -1654 593593 -1418 593829
rect -1974 593273 -1738 593509
rect -1654 593273 -1418 593509
rect 19952 593593 20188 593829
rect 19952 593273 20188 593509
rect 25882 593593 26118 593829
rect 25882 593273 26118 593509
rect 31813 593593 32049 593829
rect 31813 593273 32049 593509
rect 47952 593593 48188 593829
rect 47952 593273 48188 593509
rect 53882 593593 54118 593829
rect 53882 593273 54118 593509
rect 59813 593593 60049 593829
rect 59813 593273 60049 593509
rect 75952 593593 76188 593829
rect 75952 593273 76188 593509
rect 81882 593593 82118 593829
rect 81882 593273 82118 593509
rect 87813 593593 88049 593829
rect 87813 593273 88049 593509
rect 103952 593593 104188 593829
rect 103952 593273 104188 593509
rect 109882 593593 110118 593829
rect 109882 593273 110118 593509
rect 115813 593593 116049 593829
rect 115813 593273 116049 593509
rect 131952 593593 132188 593829
rect 131952 593273 132188 593509
rect 137882 593593 138118 593829
rect 137882 593273 138118 593509
rect 143813 593593 144049 593829
rect 143813 593273 144049 593509
rect 159952 593593 160188 593829
rect 159952 593273 160188 593509
rect 165882 593593 166118 593829
rect 165882 593273 166118 593509
rect 171813 593593 172049 593829
rect 171813 593273 172049 593509
rect 187952 593593 188188 593829
rect 187952 593273 188188 593509
rect 193882 593593 194118 593829
rect 193882 593273 194118 593509
rect 199813 593593 200049 593829
rect 199813 593273 200049 593509
rect 215952 593593 216188 593829
rect 215952 593273 216188 593509
rect 221882 593593 222118 593829
rect 221882 593273 222118 593509
rect 227813 593593 228049 593829
rect 227813 593273 228049 593509
rect 243952 593593 244188 593829
rect 243952 593273 244188 593509
rect 249882 593593 250118 593829
rect 249882 593273 250118 593509
rect 255813 593593 256049 593829
rect 255813 593273 256049 593509
rect 271952 593593 272188 593829
rect 271952 593273 272188 593509
rect 277882 593593 278118 593829
rect 277882 593273 278118 593509
rect 283813 593593 284049 593829
rect 283813 593273 284049 593509
rect 299952 593593 300188 593829
rect 299952 593273 300188 593509
rect 305882 593593 306118 593829
rect 305882 593273 306118 593509
rect 311813 593593 312049 593829
rect 311813 593273 312049 593509
rect 327952 593593 328188 593829
rect 327952 593273 328188 593509
rect 333882 593593 334118 593829
rect 333882 593273 334118 593509
rect 339813 593593 340049 593829
rect 339813 593273 340049 593509
rect 355952 593593 356188 593829
rect 355952 593273 356188 593509
rect 361882 593593 362118 593829
rect 361882 593273 362118 593509
rect 367813 593593 368049 593829
rect 367813 593273 368049 593509
rect 383952 593593 384188 593829
rect 383952 593273 384188 593509
rect 389882 593593 390118 593829
rect 389882 593273 390118 593509
rect 395813 593593 396049 593829
rect 395813 593273 396049 593509
rect 411952 593593 412188 593829
rect 411952 593273 412188 593509
rect 417882 593593 418118 593829
rect 417882 593273 418118 593509
rect 423813 593593 424049 593829
rect 423813 593273 424049 593509
rect 439952 593593 440188 593829
rect 439952 593273 440188 593509
rect 445882 593593 446118 593829
rect 445882 593273 446118 593509
rect 451813 593593 452049 593829
rect 451813 593273 452049 593509
rect 467952 593593 468188 593829
rect 467952 593273 468188 593509
rect 473882 593593 474118 593829
rect 473882 593273 474118 593509
rect 479813 593593 480049 593829
rect 479813 593273 480049 593509
rect 495952 593593 496188 593829
rect 495952 593273 496188 593509
rect 501882 593593 502118 593829
rect 501882 593273 502118 593509
rect 507813 593593 508049 593829
rect 507813 593273 508049 593509
rect 523952 593593 524188 593829
rect 523952 593273 524188 593509
rect 529882 593593 530118 593829
rect 529882 593273 530118 593509
rect 535813 593593 536049 593829
rect 535813 593273 536049 593509
rect 551952 593593 552188 593829
rect 551952 593273 552188 593509
rect 557882 593593 558118 593829
rect 557882 593273 558118 593509
rect 563813 593593 564049 593829
rect 563813 593273 564049 593509
rect 573526 593593 573762 593829
rect 573846 593593 574082 593829
rect 573526 593273 573762 593509
rect 573846 593273 574082 593509
rect 22916 590218 23152 590454
rect 22916 589898 23152 590134
rect 28847 590218 29083 590454
rect 28847 589898 29083 590134
rect 50916 590218 51152 590454
rect 50916 589898 51152 590134
rect 56847 590218 57083 590454
rect 56847 589898 57083 590134
rect 78916 590218 79152 590454
rect 78916 589898 79152 590134
rect 84847 590218 85083 590454
rect 84847 589898 85083 590134
rect 106916 590218 107152 590454
rect 106916 589898 107152 590134
rect 112847 590218 113083 590454
rect 112847 589898 113083 590134
rect 134916 590218 135152 590454
rect 134916 589898 135152 590134
rect 140847 590218 141083 590454
rect 140847 589898 141083 590134
rect 162916 590218 163152 590454
rect 162916 589898 163152 590134
rect 168847 590218 169083 590454
rect 168847 589898 169083 590134
rect 190916 590218 191152 590454
rect 190916 589898 191152 590134
rect 196847 590218 197083 590454
rect 196847 589898 197083 590134
rect 218916 590218 219152 590454
rect 218916 589898 219152 590134
rect 224847 590218 225083 590454
rect 224847 589898 225083 590134
rect 246916 590218 247152 590454
rect 246916 589898 247152 590134
rect 252847 590218 253083 590454
rect 252847 589898 253083 590134
rect 274916 590218 275152 590454
rect 274916 589898 275152 590134
rect 280847 590218 281083 590454
rect 280847 589898 281083 590134
rect 302916 590218 303152 590454
rect 302916 589898 303152 590134
rect 308847 590218 309083 590454
rect 308847 589898 309083 590134
rect 330916 590218 331152 590454
rect 330916 589898 331152 590134
rect 336847 590218 337083 590454
rect 336847 589898 337083 590134
rect 358916 590218 359152 590454
rect 358916 589898 359152 590134
rect 364847 590218 365083 590454
rect 364847 589898 365083 590134
rect 386916 590218 387152 590454
rect 386916 589898 387152 590134
rect 392847 590218 393083 590454
rect 392847 589898 393083 590134
rect 414916 590218 415152 590454
rect 414916 589898 415152 590134
rect 420847 590218 421083 590454
rect 420847 589898 421083 590134
rect 442916 590218 443152 590454
rect 442916 589898 443152 590134
rect 448847 590218 449083 590454
rect 448847 589898 449083 590134
rect 470916 590218 471152 590454
rect 470916 589898 471152 590134
rect 476847 590218 477083 590454
rect 476847 589898 477083 590134
rect 498916 590218 499152 590454
rect 498916 589898 499152 590134
rect 504847 590218 505083 590454
rect 504847 589898 505083 590134
rect 526916 590218 527152 590454
rect 526916 589898 527152 590134
rect 532847 590218 533083 590454
rect 532847 589898 533083 590134
rect 554916 590218 555152 590454
rect 554916 589898 555152 590134
rect 560847 590218 561083 590454
rect 560847 589898 561083 590134
rect -1974 566593 -1738 566829
rect -1654 566593 -1418 566829
rect -1974 566273 -1738 566509
rect -1654 566273 -1418 566509
rect 19952 566593 20188 566829
rect 19952 566273 20188 566509
rect 25882 566593 26118 566829
rect 25882 566273 26118 566509
rect 31813 566593 32049 566829
rect 31813 566273 32049 566509
rect 47952 566593 48188 566829
rect 47952 566273 48188 566509
rect 53882 566593 54118 566829
rect 53882 566273 54118 566509
rect 59813 566593 60049 566829
rect 59813 566273 60049 566509
rect 75952 566593 76188 566829
rect 75952 566273 76188 566509
rect 81882 566593 82118 566829
rect 81882 566273 82118 566509
rect 87813 566593 88049 566829
rect 87813 566273 88049 566509
rect 103952 566593 104188 566829
rect 103952 566273 104188 566509
rect 109882 566593 110118 566829
rect 109882 566273 110118 566509
rect 115813 566593 116049 566829
rect 115813 566273 116049 566509
rect 131952 566593 132188 566829
rect 131952 566273 132188 566509
rect 137882 566593 138118 566829
rect 137882 566273 138118 566509
rect 143813 566593 144049 566829
rect 143813 566273 144049 566509
rect 159952 566593 160188 566829
rect 159952 566273 160188 566509
rect 165882 566593 166118 566829
rect 165882 566273 166118 566509
rect 171813 566593 172049 566829
rect 171813 566273 172049 566509
rect 187952 566593 188188 566829
rect 187952 566273 188188 566509
rect 193882 566593 194118 566829
rect 193882 566273 194118 566509
rect 199813 566593 200049 566829
rect 199813 566273 200049 566509
rect 215952 566593 216188 566829
rect 215952 566273 216188 566509
rect 221882 566593 222118 566829
rect 221882 566273 222118 566509
rect 227813 566593 228049 566829
rect 227813 566273 228049 566509
rect 243952 566593 244188 566829
rect 243952 566273 244188 566509
rect 249882 566593 250118 566829
rect 249882 566273 250118 566509
rect 255813 566593 256049 566829
rect 255813 566273 256049 566509
rect 271952 566593 272188 566829
rect 271952 566273 272188 566509
rect 277882 566593 278118 566829
rect 277882 566273 278118 566509
rect 283813 566593 284049 566829
rect 283813 566273 284049 566509
rect 299952 566593 300188 566829
rect 299952 566273 300188 566509
rect 305882 566593 306118 566829
rect 305882 566273 306118 566509
rect 311813 566593 312049 566829
rect 311813 566273 312049 566509
rect 327952 566593 328188 566829
rect 327952 566273 328188 566509
rect 333882 566593 334118 566829
rect 333882 566273 334118 566509
rect 339813 566593 340049 566829
rect 339813 566273 340049 566509
rect 355952 566593 356188 566829
rect 355952 566273 356188 566509
rect 361882 566593 362118 566829
rect 361882 566273 362118 566509
rect 367813 566593 368049 566829
rect 367813 566273 368049 566509
rect 383952 566593 384188 566829
rect 383952 566273 384188 566509
rect 389882 566593 390118 566829
rect 389882 566273 390118 566509
rect 395813 566593 396049 566829
rect 395813 566273 396049 566509
rect 411952 566593 412188 566829
rect 411952 566273 412188 566509
rect 417882 566593 418118 566829
rect 417882 566273 418118 566509
rect 423813 566593 424049 566829
rect 423813 566273 424049 566509
rect 439952 566593 440188 566829
rect 439952 566273 440188 566509
rect 445882 566593 446118 566829
rect 445882 566273 446118 566509
rect 451813 566593 452049 566829
rect 451813 566273 452049 566509
rect 467952 566593 468188 566829
rect 467952 566273 468188 566509
rect 473882 566593 474118 566829
rect 473882 566273 474118 566509
rect 479813 566593 480049 566829
rect 479813 566273 480049 566509
rect 495952 566593 496188 566829
rect 495952 566273 496188 566509
rect 501882 566593 502118 566829
rect 501882 566273 502118 566509
rect 507813 566593 508049 566829
rect 507813 566273 508049 566509
rect 523952 566593 524188 566829
rect 523952 566273 524188 566509
rect 529882 566593 530118 566829
rect 529882 566273 530118 566509
rect 535813 566593 536049 566829
rect 535813 566273 536049 566509
rect 551952 566593 552188 566829
rect 551952 566273 552188 566509
rect 557882 566593 558118 566829
rect 557882 566273 558118 566509
rect 563813 566593 564049 566829
rect 563813 566273 564049 566509
rect 573526 566593 573762 566829
rect 573846 566593 574082 566829
rect 573526 566273 573762 566509
rect 573846 566273 574082 566509
rect 22916 563218 23152 563454
rect 22916 562898 23152 563134
rect 28847 563218 29083 563454
rect 28847 562898 29083 563134
rect 50916 563218 51152 563454
rect 50916 562898 51152 563134
rect 56847 563218 57083 563454
rect 56847 562898 57083 563134
rect 78916 563218 79152 563454
rect 78916 562898 79152 563134
rect 84847 563218 85083 563454
rect 84847 562898 85083 563134
rect 106916 563218 107152 563454
rect 106916 562898 107152 563134
rect 112847 563218 113083 563454
rect 112847 562898 113083 563134
rect 134916 563218 135152 563454
rect 134916 562898 135152 563134
rect 140847 563218 141083 563454
rect 140847 562898 141083 563134
rect 162916 563218 163152 563454
rect 162916 562898 163152 563134
rect 168847 563218 169083 563454
rect 168847 562898 169083 563134
rect 190916 563218 191152 563454
rect 190916 562898 191152 563134
rect 196847 563218 197083 563454
rect 196847 562898 197083 563134
rect 218916 563218 219152 563454
rect 218916 562898 219152 563134
rect 224847 563218 225083 563454
rect 224847 562898 225083 563134
rect 246916 563218 247152 563454
rect 246916 562898 247152 563134
rect 252847 563218 253083 563454
rect 252847 562898 253083 563134
rect 274916 563218 275152 563454
rect 274916 562898 275152 563134
rect 280847 563218 281083 563454
rect 280847 562898 281083 563134
rect 302916 563218 303152 563454
rect 302916 562898 303152 563134
rect 308847 563218 309083 563454
rect 308847 562898 309083 563134
rect 330916 563218 331152 563454
rect 330916 562898 331152 563134
rect 336847 563218 337083 563454
rect 336847 562898 337083 563134
rect 358916 563218 359152 563454
rect 358916 562898 359152 563134
rect 364847 563218 365083 563454
rect 364847 562898 365083 563134
rect 386916 563218 387152 563454
rect 386916 562898 387152 563134
rect 392847 563218 393083 563454
rect 392847 562898 393083 563134
rect 414916 563218 415152 563454
rect 414916 562898 415152 563134
rect 420847 563218 421083 563454
rect 420847 562898 421083 563134
rect 442916 563218 443152 563454
rect 442916 562898 443152 563134
rect 448847 563218 449083 563454
rect 448847 562898 449083 563134
rect 470916 563218 471152 563454
rect 470916 562898 471152 563134
rect 476847 563218 477083 563454
rect 476847 562898 477083 563134
rect 498916 563218 499152 563454
rect 498916 562898 499152 563134
rect 504847 563218 505083 563454
rect 504847 562898 505083 563134
rect 526916 563218 527152 563454
rect 526916 562898 527152 563134
rect 532847 563218 533083 563454
rect 532847 562898 533083 563134
rect 554916 563218 555152 563454
rect 554916 562898 555152 563134
rect 560847 563218 561083 563454
rect 560847 562898 561083 563134
rect -1974 539593 -1738 539829
rect -1654 539593 -1418 539829
rect -1974 539273 -1738 539509
rect -1654 539273 -1418 539509
rect 19952 539593 20188 539829
rect 19952 539273 20188 539509
rect 25882 539593 26118 539829
rect 25882 539273 26118 539509
rect 31813 539593 32049 539829
rect 31813 539273 32049 539509
rect 47952 539593 48188 539829
rect 47952 539273 48188 539509
rect 53882 539593 54118 539829
rect 53882 539273 54118 539509
rect 59813 539593 60049 539829
rect 59813 539273 60049 539509
rect 75952 539593 76188 539829
rect 75952 539273 76188 539509
rect 81882 539593 82118 539829
rect 81882 539273 82118 539509
rect 87813 539593 88049 539829
rect 87813 539273 88049 539509
rect 103952 539593 104188 539829
rect 103952 539273 104188 539509
rect 109882 539593 110118 539829
rect 109882 539273 110118 539509
rect 115813 539593 116049 539829
rect 115813 539273 116049 539509
rect 131952 539593 132188 539829
rect 131952 539273 132188 539509
rect 137882 539593 138118 539829
rect 137882 539273 138118 539509
rect 143813 539593 144049 539829
rect 143813 539273 144049 539509
rect 159952 539593 160188 539829
rect 159952 539273 160188 539509
rect 165882 539593 166118 539829
rect 165882 539273 166118 539509
rect 171813 539593 172049 539829
rect 171813 539273 172049 539509
rect 187952 539593 188188 539829
rect 187952 539273 188188 539509
rect 193882 539593 194118 539829
rect 193882 539273 194118 539509
rect 199813 539593 200049 539829
rect 199813 539273 200049 539509
rect 215952 539593 216188 539829
rect 215952 539273 216188 539509
rect 221882 539593 222118 539829
rect 221882 539273 222118 539509
rect 227813 539593 228049 539829
rect 227813 539273 228049 539509
rect 243952 539593 244188 539829
rect 243952 539273 244188 539509
rect 249882 539593 250118 539829
rect 249882 539273 250118 539509
rect 255813 539593 256049 539829
rect 255813 539273 256049 539509
rect 271952 539593 272188 539829
rect 271952 539273 272188 539509
rect 277882 539593 278118 539829
rect 277882 539273 278118 539509
rect 283813 539593 284049 539829
rect 283813 539273 284049 539509
rect 299952 539593 300188 539829
rect 299952 539273 300188 539509
rect 305882 539593 306118 539829
rect 305882 539273 306118 539509
rect 311813 539593 312049 539829
rect 311813 539273 312049 539509
rect 327952 539593 328188 539829
rect 327952 539273 328188 539509
rect 333882 539593 334118 539829
rect 333882 539273 334118 539509
rect 339813 539593 340049 539829
rect 339813 539273 340049 539509
rect 355952 539593 356188 539829
rect 355952 539273 356188 539509
rect 361882 539593 362118 539829
rect 361882 539273 362118 539509
rect 367813 539593 368049 539829
rect 367813 539273 368049 539509
rect 383952 539593 384188 539829
rect 383952 539273 384188 539509
rect 389882 539593 390118 539829
rect 389882 539273 390118 539509
rect 395813 539593 396049 539829
rect 395813 539273 396049 539509
rect 411952 539593 412188 539829
rect 411952 539273 412188 539509
rect 417882 539593 418118 539829
rect 417882 539273 418118 539509
rect 423813 539593 424049 539829
rect 423813 539273 424049 539509
rect 439952 539593 440188 539829
rect 439952 539273 440188 539509
rect 445882 539593 446118 539829
rect 445882 539273 446118 539509
rect 451813 539593 452049 539829
rect 451813 539273 452049 539509
rect 467952 539593 468188 539829
rect 467952 539273 468188 539509
rect 473882 539593 474118 539829
rect 473882 539273 474118 539509
rect 479813 539593 480049 539829
rect 479813 539273 480049 539509
rect 495952 539593 496188 539829
rect 495952 539273 496188 539509
rect 501882 539593 502118 539829
rect 501882 539273 502118 539509
rect 507813 539593 508049 539829
rect 507813 539273 508049 539509
rect 523952 539593 524188 539829
rect 523952 539273 524188 539509
rect 529882 539593 530118 539829
rect 529882 539273 530118 539509
rect 535813 539593 536049 539829
rect 535813 539273 536049 539509
rect 551952 539593 552188 539829
rect 551952 539273 552188 539509
rect 557882 539593 558118 539829
rect 557882 539273 558118 539509
rect 563813 539593 564049 539829
rect 563813 539273 564049 539509
rect 573526 539593 573762 539829
rect 573846 539593 574082 539829
rect 573526 539273 573762 539509
rect 573846 539273 574082 539509
rect 22916 536218 23152 536454
rect 22916 535898 23152 536134
rect 28847 536218 29083 536454
rect 28847 535898 29083 536134
rect 50916 536218 51152 536454
rect 50916 535898 51152 536134
rect 56847 536218 57083 536454
rect 56847 535898 57083 536134
rect 78916 536218 79152 536454
rect 78916 535898 79152 536134
rect 84847 536218 85083 536454
rect 84847 535898 85083 536134
rect 106916 536218 107152 536454
rect 106916 535898 107152 536134
rect 112847 536218 113083 536454
rect 112847 535898 113083 536134
rect 134916 536218 135152 536454
rect 134916 535898 135152 536134
rect 140847 536218 141083 536454
rect 140847 535898 141083 536134
rect 162916 536218 163152 536454
rect 162916 535898 163152 536134
rect 168847 536218 169083 536454
rect 168847 535898 169083 536134
rect 190916 536218 191152 536454
rect 190916 535898 191152 536134
rect 196847 536218 197083 536454
rect 196847 535898 197083 536134
rect 218916 536218 219152 536454
rect 218916 535898 219152 536134
rect 224847 536218 225083 536454
rect 224847 535898 225083 536134
rect 246916 536218 247152 536454
rect 246916 535898 247152 536134
rect 252847 536218 253083 536454
rect 252847 535898 253083 536134
rect 274916 536218 275152 536454
rect 274916 535898 275152 536134
rect 280847 536218 281083 536454
rect 280847 535898 281083 536134
rect 302916 536218 303152 536454
rect 302916 535898 303152 536134
rect 308847 536218 309083 536454
rect 308847 535898 309083 536134
rect 330916 536218 331152 536454
rect 330916 535898 331152 536134
rect 336847 536218 337083 536454
rect 336847 535898 337083 536134
rect 358916 536218 359152 536454
rect 358916 535898 359152 536134
rect 364847 536218 365083 536454
rect 364847 535898 365083 536134
rect 386916 536218 387152 536454
rect 386916 535898 387152 536134
rect 392847 536218 393083 536454
rect 392847 535898 393083 536134
rect 414916 536218 415152 536454
rect 414916 535898 415152 536134
rect 420847 536218 421083 536454
rect 420847 535898 421083 536134
rect 442916 536218 443152 536454
rect 442916 535898 443152 536134
rect 448847 536218 449083 536454
rect 448847 535898 449083 536134
rect 470916 536218 471152 536454
rect 470916 535898 471152 536134
rect 476847 536218 477083 536454
rect 476847 535898 477083 536134
rect 498916 536218 499152 536454
rect 498916 535898 499152 536134
rect 504847 536218 505083 536454
rect 504847 535898 505083 536134
rect 526916 536218 527152 536454
rect 526916 535898 527152 536134
rect 532847 536218 533083 536454
rect 532847 535898 533083 536134
rect 554916 536218 555152 536454
rect 554916 535898 555152 536134
rect 560847 536218 561083 536454
rect 560847 535898 561083 536134
rect -1974 512593 -1738 512829
rect -1654 512593 -1418 512829
rect -1974 512273 -1738 512509
rect -1654 512273 -1418 512509
rect 19952 512593 20188 512829
rect 19952 512273 20188 512509
rect 25882 512593 26118 512829
rect 25882 512273 26118 512509
rect 31813 512593 32049 512829
rect 31813 512273 32049 512509
rect 47952 512593 48188 512829
rect 47952 512273 48188 512509
rect 53882 512593 54118 512829
rect 53882 512273 54118 512509
rect 59813 512593 60049 512829
rect 59813 512273 60049 512509
rect 75952 512593 76188 512829
rect 75952 512273 76188 512509
rect 81882 512593 82118 512829
rect 81882 512273 82118 512509
rect 87813 512593 88049 512829
rect 87813 512273 88049 512509
rect 103952 512593 104188 512829
rect 103952 512273 104188 512509
rect 109882 512593 110118 512829
rect 109882 512273 110118 512509
rect 115813 512593 116049 512829
rect 115813 512273 116049 512509
rect 131952 512593 132188 512829
rect 131952 512273 132188 512509
rect 137882 512593 138118 512829
rect 137882 512273 138118 512509
rect 143813 512593 144049 512829
rect 143813 512273 144049 512509
rect 159952 512593 160188 512829
rect 159952 512273 160188 512509
rect 165882 512593 166118 512829
rect 165882 512273 166118 512509
rect 171813 512593 172049 512829
rect 171813 512273 172049 512509
rect 187952 512593 188188 512829
rect 187952 512273 188188 512509
rect 193882 512593 194118 512829
rect 193882 512273 194118 512509
rect 199813 512593 200049 512829
rect 199813 512273 200049 512509
rect 215952 512593 216188 512829
rect 215952 512273 216188 512509
rect 221882 512593 222118 512829
rect 221882 512273 222118 512509
rect 227813 512593 228049 512829
rect 227813 512273 228049 512509
rect 243952 512593 244188 512829
rect 243952 512273 244188 512509
rect 249882 512593 250118 512829
rect 249882 512273 250118 512509
rect 255813 512593 256049 512829
rect 255813 512273 256049 512509
rect 271952 512593 272188 512829
rect 271952 512273 272188 512509
rect 277882 512593 278118 512829
rect 277882 512273 278118 512509
rect 283813 512593 284049 512829
rect 283813 512273 284049 512509
rect 299952 512593 300188 512829
rect 299952 512273 300188 512509
rect 305882 512593 306118 512829
rect 305882 512273 306118 512509
rect 311813 512593 312049 512829
rect 311813 512273 312049 512509
rect 327952 512593 328188 512829
rect 327952 512273 328188 512509
rect 333882 512593 334118 512829
rect 333882 512273 334118 512509
rect 339813 512593 340049 512829
rect 339813 512273 340049 512509
rect 355952 512593 356188 512829
rect 355952 512273 356188 512509
rect 361882 512593 362118 512829
rect 361882 512273 362118 512509
rect 367813 512593 368049 512829
rect 367813 512273 368049 512509
rect 383952 512593 384188 512829
rect 383952 512273 384188 512509
rect 389882 512593 390118 512829
rect 389882 512273 390118 512509
rect 395813 512593 396049 512829
rect 395813 512273 396049 512509
rect 411952 512593 412188 512829
rect 411952 512273 412188 512509
rect 417882 512593 418118 512829
rect 417882 512273 418118 512509
rect 423813 512593 424049 512829
rect 423813 512273 424049 512509
rect 439952 512593 440188 512829
rect 439952 512273 440188 512509
rect 445882 512593 446118 512829
rect 445882 512273 446118 512509
rect 451813 512593 452049 512829
rect 451813 512273 452049 512509
rect 467952 512593 468188 512829
rect 467952 512273 468188 512509
rect 473882 512593 474118 512829
rect 473882 512273 474118 512509
rect 479813 512593 480049 512829
rect 479813 512273 480049 512509
rect 495952 512593 496188 512829
rect 495952 512273 496188 512509
rect 501882 512593 502118 512829
rect 501882 512273 502118 512509
rect 507813 512593 508049 512829
rect 507813 512273 508049 512509
rect 523952 512593 524188 512829
rect 523952 512273 524188 512509
rect 529882 512593 530118 512829
rect 529882 512273 530118 512509
rect 535813 512593 536049 512829
rect 535813 512273 536049 512509
rect 551952 512593 552188 512829
rect 551952 512273 552188 512509
rect 557882 512593 558118 512829
rect 557882 512273 558118 512509
rect 563813 512593 564049 512829
rect 563813 512273 564049 512509
rect 573526 512593 573762 512829
rect 573846 512593 574082 512829
rect 573526 512273 573762 512509
rect 573846 512273 574082 512509
rect 22916 509218 23152 509454
rect 22916 508898 23152 509134
rect 28847 509218 29083 509454
rect 28847 508898 29083 509134
rect 50916 509218 51152 509454
rect 50916 508898 51152 509134
rect 56847 509218 57083 509454
rect 56847 508898 57083 509134
rect 78916 509218 79152 509454
rect 78916 508898 79152 509134
rect 84847 509218 85083 509454
rect 84847 508898 85083 509134
rect 106916 509218 107152 509454
rect 106916 508898 107152 509134
rect 112847 509218 113083 509454
rect 112847 508898 113083 509134
rect 134916 509218 135152 509454
rect 134916 508898 135152 509134
rect 140847 509218 141083 509454
rect 140847 508898 141083 509134
rect 162916 509218 163152 509454
rect 162916 508898 163152 509134
rect 168847 509218 169083 509454
rect 168847 508898 169083 509134
rect 190916 509218 191152 509454
rect 190916 508898 191152 509134
rect 196847 509218 197083 509454
rect 196847 508898 197083 509134
rect 218916 509218 219152 509454
rect 218916 508898 219152 509134
rect 224847 509218 225083 509454
rect 224847 508898 225083 509134
rect 246916 509218 247152 509454
rect 246916 508898 247152 509134
rect 252847 509218 253083 509454
rect 252847 508898 253083 509134
rect 274916 509218 275152 509454
rect 274916 508898 275152 509134
rect 280847 509218 281083 509454
rect 280847 508898 281083 509134
rect 302916 509218 303152 509454
rect 302916 508898 303152 509134
rect 308847 509218 309083 509454
rect 308847 508898 309083 509134
rect 330916 509218 331152 509454
rect 330916 508898 331152 509134
rect 336847 509218 337083 509454
rect 336847 508898 337083 509134
rect 358916 509218 359152 509454
rect 358916 508898 359152 509134
rect 364847 509218 365083 509454
rect 364847 508898 365083 509134
rect 386916 509218 387152 509454
rect 386916 508898 387152 509134
rect 392847 509218 393083 509454
rect 392847 508898 393083 509134
rect 414916 509218 415152 509454
rect 414916 508898 415152 509134
rect 420847 509218 421083 509454
rect 420847 508898 421083 509134
rect 442916 509218 443152 509454
rect 442916 508898 443152 509134
rect 448847 509218 449083 509454
rect 448847 508898 449083 509134
rect 470916 509218 471152 509454
rect 470916 508898 471152 509134
rect 476847 509218 477083 509454
rect 476847 508898 477083 509134
rect 498916 509218 499152 509454
rect 498916 508898 499152 509134
rect 504847 509218 505083 509454
rect 504847 508898 505083 509134
rect 526916 509218 527152 509454
rect 526916 508898 527152 509134
rect 532847 509218 533083 509454
rect 532847 508898 533083 509134
rect 554916 509218 555152 509454
rect 554916 508898 555152 509134
rect 560847 509218 561083 509454
rect 560847 508898 561083 509134
rect -1974 485593 -1738 485829
rect -1654 485593 -1418 485829
rect -1974 485273 -1738 485509
rect -1654 485273 -1418 485509
rect 19952 485593 20188 485829
rect 19952 485273 20188 485509
rect 25882 485593 26118 485829
rect 25882 485273 26118 485509
rect 31813 485593 32049 485829
rect 31813 485273 32049 485509
rect 47952 485593 48188 485829
rect 47952 485273 48188 485509
rect 53882 485593 54118 485829
rect 53882 485273 54118 485509
rect 59813 485593 60049 485829
rect 59813 485273 60049 485509
rect 75952 485593 76188 485829
rect 75952 485273 76188 485509
rect 81882 485593 82118 485829
rect 81882 485273 82118 485509
rect 87813 485593 88049 485829
rect 87813 485273 88049 485509
rect 103952 485593 104188 485829
rect 103952 485273 104188 485509
rect 109882 485593 110118 485829
rect 109882 485273 110118 485509
rect 115813 485593 116049 485829
rect 115813 485273 116049 485509
rect 131952 485593 132188 485829
rect 131952 485273 132188 485509
rect 137882 485593 138118 485829
rect 137882 485273 138118 485509
rect 143813 485593 144049 485829
rect 143813 485273 144049 485509
rect 159952 485593 160188 485829
rect 159952 485273 160188 485509
rect 165882 485593 166118 485829
rect 165882 485273 166118 485509
rect 171813 485593 172049 485829
rect 171813 485273 172049 485509
rect 187952 485593 188188 485829
rect 187952 485273 188188 485509
rect 193882 485593 194118 485829
rect 193882 485273 194118 485509
rect 199813 485593 200049 485829
rect 199813 485273 200049 485509
rect 215952 485593 216188 485829
rect 215952 485273 216188 485509
rect 221882 485593 222118 485829
rect 221882 485273 222118 485509
rect 227813 485593 228049 485829
rect 227813 485273 228049 485509
rect 243952 485593 244188 485829
rect 243952 485273 244188 485509
rect 249882 485593 250118 485829
rect 249882 485273 250118 485509
rect 255813 485593 256049 485829
rect 255813 485273 256049 485509
rect 271952 485593 272188 485829
rect 271952 485273 272188 485509
rect 277882 485593 278118 485829
rect 277882 485273 278118 485509
rect 283813 485593 284049 485829
rect 283813 485273 284049 485509
rect 299952 485593 300188 485829
rect 299952 485273 300188 485509
rect 305882 485593 306118 485829
rect 305882 485273 306118 485509
rect 311813 485593 312049 485829
rect 311813 485273 312049 485509
rect 327952 485593 328188 485829
rect 327952 485273 328188 485509
rect 333882 485593 334118 485829
rect 333882 485273 334118 485509
rect 339813 485593 340049 485829
rect 339813 485273 340049 485509
rect 355952 485593 356188 485829
rect 355952 485273 356188 485509
rect 361882 485593 362118 485829
rect 361882 485273 362118 485509
rect 367813 485593 368049 485829
rect 367813 485273 368049 485509
rect 383952 485593 384188 485829
rect 383952 485273 384188 485509
rect 389882 485593 390118 485829
rect 389882 485273 390118 485509
rect 395813 485593 396049 485829
rect 395813 485273 396049 485509
rect 411952 485593 412188 485829
rect 411952 485273 412188 485509
rect 417882 485593 418118 485829
rect 417882 485273 418118 485509
rect 423813 485593 424049 485829
rect 423813 485273 424049 485509
rect 439952 485593 440188 485829
rect 439952 485273 440188 485509
rect 445882 485593 446118 485829
rect 445882 485273 446118 485509
rect 451813 485593 452049 485829
rect 451813 485273 452049 485509
rect 467952 485593 468188 485829
rect 467952 485273 468188 485509
rect 473882 485593 474118 485829
rect 473882 485273 474118 485509
rect 479813 485593 480049 485829
rect 479813 485273 480049 485509
rect 495952 485593 496188 485829
rect 495952 485273 496188 485509
rect 501882 485593 502118 485829
rect 501882 485273 502118 485509
rect 507813 485593 508049 485829
rect 507813 485273 508049 485509
rect 523952 485593 524188 485829
rect 523952 485273 524188 485509
rect 529882 485593 530118 485829
rect 529882 485273 530118 485509
rect 535813 485593 536049 485829
rect 535813 485273 536049 485509
rect 551952 485593 552188 485829
rect 551952 485273 552188 485509
rect 557882 485593 558118 485829
rect 557882 485273 558118 485509
rect 563813 485593 564049 485829
rect 563813 485273 564049 485509
rect 573526 485593 573762 485829
rect 573846 485593 574082 485829
rect 573526 485273 573762 485509
rect 573846 485273 574082 485509
rect 22916 482218 23152 482454
rect 22916 481898 23152 482134
rect 28847 482218 29083 482454
rect 28847 481898 29083 482134
rect 50916 482218 51152 482454
rect 50916 481898 51152 482134
rect 56847 482218 57083 482454
rect 56847 481898 57083 482134
rect 78916 482218 79152 482454
rect 78916 481898 79152 482134
rect 84847 482218 85083 482454
rect 84847 481898 85083 482134
rect 106916 482218 107152 482454
rect 106916 481898 107152 482134
rect 112847 482218 113083 482454
rect 112847 481898 113083 482134
rect 134916 482218 135152 482454
rect 134916 481898 135152 482134
rect 140847 482218 141083 482454
rect 140847 481898 141083 482134
rect 162916 482218 163152 482454
rect 162916 481898 163152 482134
rect 168847 482218 169083 482454
rect 168847 481898 169083 482134
rect 190916 482218 191152 482454
rect 190916 481898 191152 482134
rect 196847 482218 197083 482454
rect 196847 481898 197083 482134
rect 218916 482218 219152 482454
rect 218916 481898 219152 482134
rect 224847 482218 225083 482454
rect 224847 481898 225083 482134
rect 246916 482218 247152 482454
rect 246916 481898 247152 482134
rect 252847 482218 253083 482454
rect 252847 481898 253083 482134
rect 274916 482218 275152 482454
rect 274916 481898 275152 482134
rect 280847 482218 281083 482454
rect 280847 481898 281083 482134
rect 302916 482218 303152 482454
rect 302916 481898 303152 482134
rect 308847 482218 309083 482454
rect 308847 481898 309083 482134
rect 330916 482218 331152 482454
rect 330916 481898 331152 482134
rect 336847 482218 337083 482454
rect 336847 481898 337083 482134
rect 358916 482218 359152 482454
rect 358916 481898 359152 482134
rect 364847 482218 365083 482454
rect 364847 481898 365083 482134
rect 386916 482218 387152 482454
rect 386916 481898 387152 482134
rect 392847 482218 393083 482454
rect 392847 481898 393083 482134
rect 414916 482218 415152 482454
rect 414916 481898 415152 482134
rect 420847 482218 421083 482454
rect 420847 481898 421083 482134
rect 442916 482218 443152 482454
rect 442916 481898 443152 482134
rect 448847 482218 449083 482454
rect 448847 481898 449083 482134
rect 470916 482218 471152 482454
rect 470916 481898 471152 482134
rect 476847 482218 477083 482454
rect 476847 481898 477083 482134
rect 498916 482218 499152 482454
rect 498916 481898 499152 482134
rect 504847 482218 505083 482454
rect 504847 481898 505083 482134
rect 526916 482218 527152 482454
rect 526916 481898 527152 482134
rect 532847 482218 533083 482454
rect 532847 481898 533083 482134
rect 554916 482218 555152 482454
rect 554916 481898 555152 482134
rect 560847 482218 561083 482454
rect 560847 481898 561083 482134
rect -1974 458593 -1738 458829
rect -1654 458593 -1418 458829
rect -1974 458273 -1738 458509
rect -1654 458273 -1418 458509
rect 19952 458593 20188 458829
rect 19952 458273 20188 458509
rect 25882 458593 26118 458829
rect 25882 458273 26118 458509
rect 31813 458593 32049 458829
rect 31813 458273 32049 458509
rect 47952 458593 48188 458829
rect 47952 458273 48188 458509
rect 53882 458593 54118 458829
rect 53882 458273 54118 458509
rect 59813 458593 60049 458829
rect 59813 458273 60049 458509
rect 75952 458593 76188 458829
rect 75952 458273 76188 458509
rect 81882 458593 82118 458829
rect 81882 458273 82118 458509
rect 87813 458593 88049 458829
rect 87813 458273 88049 458509
rect 103952 458593 104188 458829
rect 103952 458273 104188 458509
rect 109882 458593 110118 458829
rect 109882 458273 110118 458509
rect 115813 458593 116049 458829
rect 115813 458273 116049 458509
rect 131952 458593 132188 458829
rect 131952 458273 132188 458509
rect 137882 458593 138118 458829
rect 137882 458273 138118 458509
rect 143813 458593 144049 458829
rect 143813 458273 144049 458509
rect 159952 458593 160188 458829
rect 159952 458273 160188 458509
rect 165882 458593 166118 458829
rect 165882 458273 166118 458509
rect 171813 458593 172049 458829
rect 171813 458273 172049 458509
rect 187952 458593 188188 458829
rect 187952 458273 188188 458509
rect 193882 458593 194118 458829
rect 193882 458273 194118 458509
rect 199813 458593 200049 458829
rect 199813 458273 200049 458509
rect 215952 458593 216188 458829
rect 215952 458273 216188 458509
rect 221882 458593 222118 458829
rect 221882 458273 222118 458509
rect 227813 458593 228049 458829
rect 227813 458273 228049 458509
rect 243952 458593 244188 458829
rect 243952 458273 244188 458509
rect 249882 458593 250118 458829
rect 249882 458273 250118 458509
rect 255813 458593 256049 458829
rect 255813 458273 256049 458509
rect 271952 458593 272188 458829
rect 271952 458273 272188 458509
rect 277882 458593 278118 458829
rect 277882 458273 278118 458509
rect 283813 458593 284049 458829
rect 283813 458273 284049 458509
rect 299952 458593 300188 458829
rect 299952 458273 300188 458509
rect 305882 458593 306118 458829
rect 305882 458273 306118 458509
rect 311813 458593 312049 458829
rect 311813 458273 312049 458509
rect 327952 458593 328188 458829
rect 327952 458273 328188 458509
rect 333882 458593 334118 458829
rect 333882 458273 334118 458509
rect 339813 458593 340049 458829
rect 339813 458273 340049 458509
rect 355952 458593 356188 458829
rect 355952 458273 356188 458509
rect 361882 458593 362118 458829
rect 361882 458273 362118 458509
rect 367813 458593 368049 458829
rect 367813 458273 368049 458509
rect 383952 458593 384188 458829
rect 383952 458273 384188 458509
rect 389882 458593 390118 458829
rect 389882 458273 390118 458509
rect 395813 458593 396049 458829
rect 395813 458273 396049 458509
rect 411952 458593 412188 458829
rect 411952 458273 412188 458509
rect 417882 458593 418118 458829
rect 417882 458273 418118 458509
rect 423813 458593 424049 458829
rect 423813 458273 424049 458509
rect 439952 458593 440188 458829
rect 439952 458273 440188 458509
rect 445882 458593 446118 458829
rect 445882 458273 446118 458509
rect 451813 458593 452049 458829
rect 451813 458273 452049 458509
rect 467952 458593 468188 458829
rect 467952 458273 468188 458509
rect 473882 458593 474118 458829
rect 473882 458273 474118 458509
rect 479813 458593 480049 458829
rect 479813 458273 480049 458509
rect 495952 458593 496188 458829
rect 495952 458273 496188 458509
rect 501882 458593 502118 458829
rect 501882 458273 502118 458509
rect 507813 458593 508049 458829
rect 507813 458273 508049 458509
rect 523952 458593 524188 458829
rect 523952 458273 524188 458509
rect 529882 458593 530118 458829
rect 529882 458273 530118 458509
rect 535813 458593 536049 458829
rect 535813 458273 536049 458509
rect 551952 458593 552188 458829
rect 551952 458273 552188 458509
rect 557882 458593 558118 458829
rect 557882 458273 558118 458509
rect 563813 458593 564049 458829
rect 563813 458273 564049 458509
rect 573526 458593 573762 458829
rect 573846 458593 574082 458829
rect 573526 458273 573762 458509
rect 573846 458273 574082 458509
rect 22916 455218 23152 455454
rect 22916 454898 23152 455134
rect 28847 455218 29083 455454
rect 28847 454898 29083 455134
rect 50916 455218 51152 455454
rect 50916 454898 51152 455134
rect 56847 455218 57083 455454
rect 56847 454898 57083 455134
rect 78916 455218 79152 455454
rect 78916 454898 79152 455134
rect 84847 455218 85083 455454
rect 84847 454898 85083 455134
rect 106916 455218 107152 455454
rect 106916 454898 107152 455134
rect 112847 455218 113083 455454
rect 112847 454898 113083 455134
rect 134916 455218 135152 455454
rect 134916 454898 135152 455134
rect 140847 455218 141083 455454
rect 140847 454898 141083 455134
rect 162916 455218 163152 455454
rect 162916 454898 163152 455134
rect 168847 455218 169083 455454
rect 168847 454898 169083 455134
rect 190916 455218 191152 455454
rect 190916 454898 191152 455134
rect 196847 455218 197083 455454
rect 196847 454898 197083 455134
rect 218916 455218 219152 455454
rect 218916 454898 219152 455134
rect 224847 455218 225083 455454
rect 224847 454898 225083 455134
rect 246916 455218 247152 455454
rect 246916 454898 247152 455134
rect 252847 455218 253083 455454
rect 252847 454898 253083 455134
rect 274916 455218 275152 455454
rect 274916 454898 275152 455134
rect 280847 455218 281083 455454
rect 280847 454898 281083 455134
rect 302916 455218 303152 455454
rect 302916 454898 303152 455134
rect 308847 455218 309083 455454
rect 308847 454898 309083 455134
rect 330916 455218 331152 455454
rect 330916 454898 331152 455134
rect 336847 455218 337083 455454
rect 336847 454898 337083 455134
rect 358916 455218 359152 455454
rect 358916 454898 359152 455134
rect 364847 455218 365083 455454
rect 364847 454898 365083 455134
rect 386916 455218 387152 455454
rect 386916 454898 387152 455134
rect 392847 455218 393083 455454
rect 392847 454898 393083 455134
rect 414916 455218 415152 455454
rect 414916 454898 415152 455134
rect 420847 455218 421083 455454
rect 420847 454898 421083 455134
rect 442916 455218 443152 455454
rect 442916 454898 443152 455134
rect 448847 455218 449083 455454
rect 448847 454898 449083 455134
rect 470916 455218 471152 455454
rect 470916 454898 471152 455134
rect 476847 455218 477083 455454
rect 476847 454898 477083 455134
rect 498916 455218 499152 455454
rect 498916 454898 499152 455134
rect 504847 455218 505083 455454
rect 504847 454898 505083 455134
rect 526916 455218 527152 455454
rect 526916 454898 527152 455134
rect 532847 455218 533083 455454
rect 532847 454898 533083 455134
rect 554916 455218 555152 455454
rect 554916 454898 555152 455134
rect 560847 455218 561083 455454
rect 560847 454898 561083 455134
rect -1974 431593 -1738 431829
rect -1654 431593 -1418 431829
rect -1974 431273 -1738 431509
rect -1654 431273 -1418 431509
rect 19952 431593 20188 431829
rect 19952 431273 20188 431509
rect 25882 431593 26118 431829
rect 25882 431273 26118 431509
rect 31813 431593 32049 431829
rect 31813 431273 32049 431509
rect 47952 431593 48188 431829
rect 47952 431273 48188 431509
rect 53882 431593 54118 431829
rect 53882 431273 54118 431509
rect 59813 431593 60049 431829
rect 59813 431273 60049 431509
rect 75952 431593 76188 431829
rect 75952 431273 76188 431509
rect 81882 431593 82118 431829
rect 81882 431273 82118 431509
rect 87813 431593 88049 431829
rect 87813 431273 88049 431509
rect 103952 431593 104188 431829
rect 103952 431273 104188 431509
rect 109882 431593 110118 431829
rect 109882 431273 110118 431509
rect 115813 431593 116049 431829
rect 115813 431273 116049 431509
rect 131952 431593 132188 431829
rect 131952 431273 132188 431509
rect 137882 431593 138118 431829
rect 137882 431273 138118 431509
rect 143813 431593 144049 431829
rect 143813 431273 144049 431509
rect 159952 431593 160188 431829
rect 159952 431273 160188 431509
rect 165882 431593 166118 431829
rect 165882 431273 166118 431509
rect 171813 431593 172049 431829
rect 171813 431273 172049 431509
rect 187952 431593 188188 431829
rect 187952 431273 188188 431509
rect 193882 431593 194118 431829
rect 193882 431273 194118 431509
rect 199813 431593 200049 431829
rect 199813 431273 200049 431509
rect 215952 431593 216188 431829
rect 215952 431273 216188 431509
rect 221882 431593 222118 431829
rect 221882 431273 222118 431509
rect 227813 431593 228049 431829
rect 227813 431273 228049 431509
rect 243952 431593 244188 431829
rect 243952 431273 244188 431509
rect 249882 431593 250118 431829
rect 249882 431273 250118 431509
rect 255813 431593 256049 431829
rect 255813 431273 256049 431509
rect 271952 431593 272188 431829
rect 271952 431273 272188 431509
rect 277882 431593 278118 431829
rect 277882 431273 278118 431509
rect 283813 431593 284049 431829
rect 283813 431273 284049 431509
rect 299952 431593 300188 431829
rect 299952 431273 300188 431509
rect 305882 431593 306118 431829
rect 305882 431273 306118 431509
rect 311813 431593 312049 431829
rect 311813 431273 312049 431509
rect 327952 431593 328188 431829
rect 327952 431273 328188 431509
rect 333882 431593 334118 431829
rect 333882 431273 334118 431509
rect 339813 431593 340049 431829
rect 339813 431273 340049 431509
rect 355952 431593 356188 431829
rect 355952 431273 356188 431509
rect 361882 431593 362118 431829
rect 361882 431273 362118 431509
rect 367813 431593 368049 431829
rect 367813 431273 368049 431509
rect 383952 431593 384188 431829
rect 383952 431273 384188 431509
rect 389882 431593 390118 431829
rect 389882 431273 390118 431509
rect 395813 431593 396049 431829
rect 395813 431273 396049 431509
rect 411952 431593 412188 431829
rect 411952 431273 412188 431509
rect 417882 431593 418118 431829
rect 417882 431273 418118 431509
rect 423813 431593 424049 431829
rect 423813 431273 424049 431509
rect 439952 431593 440188 431829
rect 439952 431273 440188 431509
rect 445882 431593 446118 431829
rect 445882 431273 446118 431509
rect 451813 431593 452049 431829
rect 451813 431273 452049 431509
rect 467952 431593 468188 431829
rect 467952 431273 468188 431509
rect 473882 431593 474118 431829
rect 473882 431273 474118 431509
rect 479813 431593 480049 431829
rect 479813 431273 480049 431509
rect 495952 431593 496188 431829
rect 495952 431273 496188 431509
rect 501882 431593 502118 431829
rect 501882 431273 502118 431509
rect 507813 431593 508049 431829
rect 507813 431273 508049 431509
rect 523952 431593 524188 431829
rect 523952 431273 524188 431509
rect 529882 431593 530118 431829
rect 529882 431273 530118 431509
rect 535813 431593 536049 431829
rect 535813 431273 536049 431509
rect 551952 431593 552188 431829
rect 551952 431273 552188 431509
rect 557882 431593 558118 431829
rect 557882 431273 558118 431509
rect 563813 431593 564049 431829
rect 563813 431273 564049 431509
rect 573526 431593 573762 431829
rect 573846 431593 574082 431829
rect 573526 431273 573762 431509
rect 573846 431273 574082 431509
rect 22916 428218 23152 428454
rect 22916 427898 23152 428134
rect 28847 428218 29083 428454
rect 28847 427898 29083 428134
rect 50916 428218 51152 428454
rect 50916 427898 51152 428134
rect 56847 428218 57083 428454
rect 56847 427898 57083 428134
rect 78916 428218 79152 428454
rect 78916 427898 79152 428134
rect 84847 428218 85083 428454
rect 84847 427898 85083 428134
rect 106916 428218 107152 428454
rect 106916 427898 107152 428134
rect 112847 428218 113083 428454
rect 112847 427898 113083 428134
rect 134916 428218 135152 428454
rect 134916 427898 135152 428134
rect 140847 428218 141083 428454
rect 140847 427898 141083 428134
rect 162916 428218 163152 428454
rect 162916 427898 163152 428134
rect 168847 428218 169083 428454
rect 168847 427898 169083 428134
rect 190916 428218 191152 428454
rect 190916 427898 191152 428134
rect 196847 428218 197083 428454
rect 196847 427898 197083 428134
rect 218916 428218 219152 428454
rect 218916 427898 219152 428134
rect 224847 428218 225083 428454
rect 224847 427898 225083 428134
rect 246916 428218 247152 428454
rect 246916 427898 247152 428134
rect 252847 428218 253083 428454
rect 252847 427898 253083 428134
rect 274916 428218 275152 428454
rect 274916 427898 275152 428134
rect 280847 428218 281083 428454
rect 280847 427898 281083 428134
rect 302916 428218 303152 428454
rect 302916 427898 303152 428134
rect 308847 428218 309083 428454
rect 308847 427898 309083 428134
rect 330916 428218 331152 428454
rect 330916 427898 331152 428134
rect 336847 428218 337083 428454
rect 336847 427898 337083 428134
rect 358916 428218 359152 428454
rect 358916 427898 359152 428134
rect 364847 428218 365083 428454
rect 364847 427898 365083 428134
rect 386916 428218 387152 428454
rect 386916 427898 387152 428134
rect 392847 428218 393083 428454
rect 392847 427898 393083 428134
rect 414916 428218 415152 428454
rect 414916 427898 415152 428134
rect 420847 428218 421083 428454
rect 420847 427898 421083 428134
rect 442916 428218 443152 428454
rect 442916 427898 443152 428134
rect 448847 428218 449083 428454
rect 448847 427898 449083 428134
rect 470916 428218 471152 428454
rect 470916 427898 471152 428134
rect 476847 428218 477083 428454
rect 476847 427898 477083 428134
rect 498916 428218 499152 428454
rect 498916 427898 499152 428134
rect 504847 428218 505083 428454
rect 504847 427898 505083 428134
rect 526916 428218 527152 428454
rect 526916 427898 527152 428134
rect 532847 428218 533083 428454
rect 532847 427898 533083 428134
rect 554916 428218 555152 428454
rect 554916 427898 555152 428134
rect 560847 428218 561083 428454
rect 560847 427898 561083 428134
rect -1974 404593 -1738 404829
rect -1654 404593 -1418 404829
rect -1974 404273 -1738 404509
rect -1654 404273 -1418 404509
rect 19952 404593 20188 404829
rect 19952 404273 20188 404509
rect 25882 404593 26118 404829
rect 25882 404273 26118 404509
rect 31813 404593 32049 404829
rect 31813 404273 32049 404509
rect 47952 404593 48188 404829
rect 47952 404273 48188 404509
rect 53882 404593 54118 404829
rect 53882 404273 54118 404509
rect 59813 404593 60049 404829
rect 59813 404273 60049 404509
rect 75952 404593 76188 404829
rect 75952 404273 76188 404509
rect 81882 404593 82118 404829
rect 81882 404273 82118 404509
rect 87813 404593 88049 404829
rect 87813 404273 88049 404509
rect 103952 404593 104188 404829
rect 103952 404273 104188 404509
rect 109882 404593 110118 404829
rect 109882 404273 110118 404509
rect 115813 404593 116049 404829
rect 115813 404273 116049 404509
rect 131952 404593 132188 404829
rect 131952 404273 132188 404509
rect 137882 404593 138118 404829
rect 137882 404273 138118 404509
rect 143813 404593 144049 404829
rect 143813 404273 144049 404509
rect 159952 404593 160188 404829
rect 159952 404273 160188 404509
rect 165882 404593 166118 404829
rect 165882 404273 166118 404509
rect 171813 404593 172049 404829
rect 171813 404273 172049 404509
rect 187952 404593 188188 404829
rect 187952 404273 188188 404509
rect 193882 404593 194118 404829
rect 193882 404273 194118 404509
rect 199813 404593 200049 404829
rect 199813 404273 200049 404509
rect 215952 404593 216188 404829
rect 215952 404273 216188 404509
rect 221882 404593 222118 404829
rect 221882 404273 222118 404509
rect 227813 404593 228049 404829
rect 227813 404273 228049 404509
rect 243952 404593 244188 404829
rect 243952 404273 244188 404509
rect 249882 404593 250118 404829
rect 249882 404273 250118 404509
rect 255813 404593 256049 404829
rect 255813 404273 256049 404509
rect 271952 404593 272188 404829
rect 271952 404273 272188 404509
rect 277882 404593 278118 404829
rect 277882 404273 278118 404509
rect 283813 404593 284049 404829
rect 283813 404273 284049 404509
rect 299952 404593 300188 404829
rect 299952 404273 300188 404509
rect 305882 404593 306118 404829
rect 305882 404273 306118 404509
rect 311813 404593 312049 404829
rect 311813 404273 312049 404509
rect 327952 404593 328188 404829
rect 327952 404273 328188 404509
rect 333882 404593 334118 404829
rect 333882 404273 334118 404509
rect 339813 404593 340049 404829
rect 339813 404273 340049 404509
rect 355952 404593 356188 404829
rect 355952 404273 356188 404509
rect 361882 404593 362118 404829
rect 361882 404273 362118 404509
rect 367813 404593 368049 404829
rect 367813 404273 368049 404509
rect 383952 404593 384188 404829
rect 383952 404273 384188 404509
rect 389882 404593 390118 404829
rect 389882 404273 390118 404509
rect 395813 404593 396049 404829
rect 395813 404273 396049 404509
rect 411952 404593 412188 404829
rect 411952 404273 412188 404509
rect 417882 404593 418118 404829
rect 417882 404273 418118 404509
rect 423813 404593 424049 404829
rect 423813 404273 424049 404509
rect 439952 404593 440188 404829
rect 439952 404273 440188 404509
rect 445882 404593 446118 404829
rect 445882 404273 446118 404509
rect 451813 404593 452049 404829
rect 451813 404273 452049 404509
rect 467952 404593 468188 404829
rect 467952 404273 468188 404509
rect 473882 404593 474118 404829
rect 473882 404273 474118 404509
rect 479813 404593 480049 404829
rect 479813 404273 480049 404509
rect 495952 404593 496188 404829
rect 495952 404273 496188 404509
rect 501882 404593 502118 404829
rect 501882 404273 502118 404509
rect 507813 404593 508049 404829
rect 507813 404273 508049 404509
rect 523952 404593 524188 404829
rect 523952 404273 524188 404509
rect 529882 404593 530118 404829
rect 529882 404273 530118 404509
rect 535813 404593 536049 404829
rect 535813 404273 536049 404509
rect 551952 404593 552188 404829
rect 551952 404273 552188 404509
rect 557882 404593 558118 404829
rect 557882 404273 558118 404509
rect 563813 404593 564049 404829
rect 563813 404273 564049 404509
rect 573526 404593 573762 404829
rect 573846 404593 574082 404829
rect 573526 404273 573762 404509
rect 573846 404273 574082 404509
rect 22916 401218 23152 401454
rect 22916 400898 23152 401134
rect 28847 401218 29083 401454
rect 28847 400898 29083 401134
rect 50916 401218 51152 401454
rect 50916 400898 51152 401134
rect 56847 401218 57083 401454
rect 56847 400898 57083 401134
rect 78916 401218 79152 401454
rect 78916 400898 79152 401134
rect 84847 401218 85083 401454
rect 84847 400898 85083 401134
rect 106916 401218 107152 401454
rect 106916 400898 107152 401134
rect 112847 401218 113083 401454
rect 112847 400898 113083 401134
rect 134916 401218 135152 401454
rect 134916 400898 135152 401134
rect 140847 401218 141083 401454
rect 140847 400898 141083 401134
rect 162916 401218 163152 401454
rect 162916 400898 163152 401134
rect 168847 401218 169083 401454
rect 168847 400898 169083 401134
rect 190916 401218 191152 401454
rect 190916 400898 191152 401134
rect 196847 401218 197083 401454
rect 196847 400898 197083 401134
rect 218916 401218 219152 401454
rect 218916 400898 219152 401134
rect 224847 401218 225083 401454
rect 224847 400898 225083 401134
rect 246916 401218 247152 401454
rect 246916 400898 247152 401134
rect 252847 401218 253083 401454
rect 252847 400898 253083 401134
rect 274916 401218 275152 401454
rect 274916 400898 275152 401134
rect 280847 401218 281083 401454
rect 280847 400898 281083 401134
rect 302916 401218 303152 401454
rect 302916 400898 303152 401134
rect 308847 401218 309083 401454
rect 308847 400898 309083 401134
rect 330916 401218 331152 401454
rect 330916 400898 331152 401134
rect 336847 401218 337083 401454
rect 336847 400898 337083 401134
rect 358916 401218 359152 401454
rect 358916 400898 359152 401134
rect 364847 401218 365083 401454
rect 364847 400898 365083 401134
rect 386916 401218 387152 401454
rect 386916 400898 387152 401134
rect 392847 401218 393083 401454
rect 392847 400898 393083 401134
rect 414916 401218 415152 401454
rect 414916 400898 415152 401134
rect 420847 401218 421083 401454
rect 420847 400898 421083 401134
rect 442916 401218 443152 401454
rect 442916 400898 443152 401134
rect 448847 401218 449083 401454
rect 448847 400898 449083 401134
rect 470916 401218 471152 401454
rect 470916 400898 471152 401134
rect 476847 401218 477083 401454
rect 476847 400898 477083 401134
rect 498916 401218 499152 401454
rect 498916 400898 499152 401134
rect 504847 401218 505083 401454
rect 504847 400898 505083 401134
rect 526916 401218 527152 401454
rect 526916 400898 527152 401134
rect 532847 401218 533083 401454
rect 532847 400898 533083 401134
rect 554916 401218 555152 401454
rect 554916 400898 555152 401134
rect 560847 401218 561083 401454
rect 560847 400898 561083 401134
rect -1974 377593 -1738 377829
rect -1654 377593 -1418 377829
rect -1974 377273 -1738 377509
rect -1654 377273 -1418 377509
rect 19952 377593 20188 377829
rect 19952 377273 20188 377509
rect 25882 377593 26118 377829
rect 25882 377273 26118 377509
rect 31813 377593 32049 377829
rect 31813 377273 32049 377509
rect 47952 377593 48188 377829
rect 47952 377273 48188 377509
rect 53882 377593 54118 377829
rect 53882 377273 54118 377509
rect 59813 377593 60049 377829
rect 59813 377273 60049 377509
rect 75952 377593 76188 377829
rect 75952 377273 76188 377509
rect 81882 377593 82118 377829
rect 81882 377273 82118 377509
rect 87813 377593 88049 377829
rect 87813 377273 88049 377509
rect 103952 377593 104188 377829
rect 103952 377273 104188 377509
rect 109882 377593 110118 377829
rect 109882 377273 110118 377509
rect 115813 377593 116049 377829
rect 115813 377273 116049 377509
rect 131952 377593 132188 377829
rect 131952 377273 132188 377509
rect 137882 377593 138118 377829
rect 137882 377273 138118 377509
rect 143813 377593 144049 377829
rect 143813 377273 144049 377509
rect 159952 377593 160188 377829
rect 159952 377273 160188 377509
rect 165882 377593 166118 377829
rect 165882 377273 166118 377509
rect 171813 377593 172049 377829
rect 171813 377273 172049 377509
rect 187952 377593 188188 377829
rect 187952 377273 188188 377509
rect 193882 377593 194118 377829
rect 193882 377273 194118 377509
rect 199813 377593 200049 377829
rect 199813 377273 200049 377509
rect 215952 377593 216188 377829
rect 215952 377273 216188 377509
rect 221882 377593 222118 377829
rect 221882 377273 222118 377509
rect 227813 377593 228049 377829
rect 227813 377273 228049 377509
rect 243952 377593 244188 377829
rect 243952 377273 244188 377509
rect 249882 377593 250118 377829
rect 249882 377273 250118 377509
rect 255813 377593 256049 377829
rect 255813 377273 256049 377509
rect 271952 377593 272188 377829
rect 271952 377273 272188 377509
rect 277882 377593 278118 377829
rect 277882 377273 278118 377509
rect 283813 377593 284049 377829
rect 283813 377273 284049 377509
rect 299952 377593 300188 377829
rect 299952 377273 300188 377509
rect 305882 377593 306118 377829
rect 305882 377273 306118 377509
rect 311813 377593 312049 377829
rect 311813 377273 312049 377509
rect 327952 377593 328188 377829
rect 327952 377273 328188 377509
rect 333882 377593 334118 377829
rect 333882 377273 334118 377509
rect 339813 377593 340049 377829
rect 339813 377273 340049 377509
rect 355952 377593 356188 377829
rect 355952 377273 356188 377509
rect 361882 377593 362118 377829
rect 361882 377273 362118 377509
rect 367813 377593 368049 377829
rect 367813 377273 368049 377509
rect 383952 377593 384188 377829
rect 383952 377273 384188 377509
rect 389882 377593 390118 377829
rect 389882 377273 390118 377509
rect 395813 377593 396049 377829
rect 395813 377273 396049 377509
rect 411952 377593 412188 377829
rect 411952 377273 412188 377509
rect 417882 377593 418118 377829
rect 417882 377273 418118 377509
rect 423813 377593 424049 377829
rect 423813 377273 424049 377509
rect 439952 377593 440188 377829
rect 439952 377273 440188 377509
rect 445882 377593 446118 377829
rect 445882 377273 446118 377509
rect 451813 377593 452049 377829
rect 451813 377273 452049 377509
rect 467952 377593 468188 377829
rect 467952 377273 468188 377509
rect 473882 377593 474118 377829
rect 473882 377273 474118 377509
rect 479813 377593 480049 377829
rect 479813 377273 480049 377509
rect 495952 377593 496188 377829
rect 495952 377273 496188 377509
rect 501882 377593 502118 377829
rect 501882 377273 502118 377509
rect 507813 377593 508049 377829
rect 507813 377273 508049 377509
rect 523952 377593 524188 377829
rect 523952 377273 524188 377509
rect 529882 377593 530118 377829
rect 529882 377273 530118 377509
rect 535813 377593 536049 377829
rect 535813 377273 536049 377509
rect 551952 377593 552188 377829
rect 551952 377273 552188 377509
rect 557882 377593 558118 377829
rect 557882 377273 558118 377509
rect 563813 377593 564049 377829
rect 563813 377273 564049 377509
rect 573526 377593 573762 377829
rect 573846 377593 574082 377829
rect 573526 377273 573762 377509
rect 573846 377273 574082 377509
rect 22916 374218 23152 374454
rect 22916 373898 23152 374134
rect 28847 374218 29083 374454
rect 28847 373898 29083 374134
rect 50916 374218 51152 374454
rect 50916 373898 51152 374134
rect 56847 374218 57083 374454
rect 56847 373898 57083 374134
rect 78916 374218 79152 374454
rect 78916 373898 79152 374134
rect 84847 374218 85083 374454
rect 84847 373898 85083 374134
rect 106916 374218 107152 374454
rect 106916 373898 107152 374134
rect 112847 374218 113083 374454
rect 112847 373898 113083 374134
rect 134916 374218 135152 374454
rect 134916 373898 135152 374134
rect 140847 374218 141083 374454
rect 140847 373898 141083 374134
rect 162916 374218 163152 374454
rect 162916 373898 163152 374134
rect 168847 374218 169083 374454
rect 168847 373898 169083 374134
rect 190916 374218 191152 374454
rect 190916 373898 191152 374134
rect 196847 374218 197083 374454
rect 196847 373898 197083 374134
rect 218916 374218 219152 374454
rect 218916 373898 219152 374134
rect 224847 374218 225083 374454
rect 224847 373898 225083 374134
rect 246916 374218 247152 374454
rect 246916 373898 247152 374134
rect 252847 374218 253083 374454
rect 252847 373898 253083 374134
rect 274916 374218 275152 374454
rect 274916 373898 275152 374134
rect 280847 374218 281083 374454
rect 280847 373898 281083 374134
rect 302916 374218 303152 374454
rect 302916 373898 303152 374134
rect 308847 374218 309083 374454
rect 308847 373898 309083 374134
rect 330916 374218 331152 374454
rect 330916 373898 331152 374134
rect 336847 374218 337083 374454
rect 336847 373898 337083 374134
rect 358916 374218 359152 374454
rect 358916 373898 359152 374134
rect 364847 374218 365083 374454
rect 364847 373898 365083 374134
rect 386916 374218 387152 374454
rect 386916 373898 387152 374134
rect 392847 374218 393083 374454
rect 392847 373898 393083 374134
rect 414916 374218 415152 374454
rect 414916 373898 415152 374134
rect 420847 374218 421083 374454
rect 420847 373898 421083 374134
rect 442916 374218 443152 374454
rect 442916 373898 443152 374134
rect 448847 374218 449083 374454
rect 448847 373898 449083 374134
rect 470916 374218 471152 374454
rect 470916 373898 471152 374134
rect 476847 374218 477083 374454
rect 476847 373898 477083 374134
rect 498916 374218 499152 374454
rect 498916 373898 499152 374134
rect 504847 374218 505083 374454
rect 504847 373898 505083 374134
rect 526916 374218 527152 374454
rect 526916 373898 527152 374134
rect 532847 374218 533083 374454
rect 532847 373898 533083 374134
rect 554916 374218 555152 374454
rect 554916 373898 555152 374134
rect 560847 374218 561083 374454
rect 560847 373898 561083 374134
rect -1974 350593 -1738 350829
rect -1654 350593 -1418 350829
rect -1974 350273 -1738 350509
rect -1654 350273 -1418 350509
rect 19952 350593 20188 350829
rect 19952 350273 20188 350509
rect 25882 350593 26118 350829
rect 25882 350273 26118 350509
rect 31813 350593 32049 350829
rect 31813 350273 32049 350509
rect 47952 350593 48188 350829
rect 47952 350273 48188 350509
rect 53882 350593 54118 350829
rect 53882 350273 54118 350509
rect 59813 350593 60049 350829
rect 59813 350273 60049 350509
rect 75952 350593 76188 350829
rect 75952 350273 76188 350509
rect 81882 350593 82118 350829
rect 81882 350273 82118 350509
rect 87813 350593 88049 350829
rect 87813 350273 88049 350509
rect 103952 350593 104188 350829
rect 103952 350273 104188 350509
rect 109882 350593 110118 350829
rect 109882 350273 110118 350509
rect 115813 350593 116049 350829
rect 115813 350273 116049 350509
rect 131952 350593 132188 350829
rect 131952 350273 132188 350509
rect 137882 350593 138118 350829
rect 137882 350273 138118 350509
rect 143813 350593 144049 350829
rect 143813 350273 144049 350509
rect 159952 350593 160188 350829
rect 159952 350273 160188 350509
rect 165882 350593 166118 350829
rect 165882 350273 166118 350509
rect 171813 350593 172049 350829
rect 171813 350273 172049 350509
rect 187952 350593 188188 350829
rect 187952 350273 188188 350509
rect 193882 350593 194118 350829
rect 193882 350273 194118 350509
rect 199813 350593 200049 350829
rect 199813 350273 200049 350509
rect 215952 350593 216188 350829
rect 215952 350273 216188 350509
rect 221882 350593 222118 350829
rect 221882 350273 222118 350509
rect 227813 350593 228049 350829
rect 227813 350273 228049 350509
rect 243952 350593 244188 350829
rect 243952 350273 244188 350509
rect 249882 350593 250118 350829
rect 249882 350273 250118 350509
rect 255813 350593 256049 350829
rect 255813 350273 256049 350509
rect 271952 350593 272188 350829
rect 271952 350273 272188 350509
rect 277882 350593 278118 350829
rect 277882 350273 278118 350509
rect 283813 350593 284049 350829
rect 283813 350273 284049 350509
rect 299952 350593 300188 350829
rect 299952 350273 300188 350509
rect 305882 350593 306118 350829
rect 305882 350273 306118 350509
rect 311813 350593 312049 350829
rect 311813 350273 312049 350509
rect 327952 350593 328188 350829
rect 327952 350273 328188 350509
rect 333882 350593 334118 350829
rect 333882 350273 334118 350509
rect 339813 350593 340049 350829
rect 339813 350273 340049 350509
rect 355952 350593 356188 350829
rect 355952 350273 356188 350509
rect 361882 350593 362118 350829
rect 361882 350273 362118 350509
rect 367813 350593 368049 350829
rect 367813 350273 368049 350509
rect 383952 350593 384188 350829
rect 383952 350273 384188 350509
rect 389882 350593 390118 350829
rect 389882 350273 390118 350509
rect 395813 350593 396049 350829
rect 395813 350273 396049 350509
rect 411952 350593 412188 350829
rect 411952 350273 412188 350509
rect 417882 350593 418118 350829
rect 417882 350273 418118 350509
rect 423813 350593 424049 350829
rect 423813 350273 424049 350509
rect 439952 350593 440188 350829
rect 439952 350273 440188 350509
rect 445882 350593 446118 350829
rect 445882 350273 446118 350509
rect 451813 350593 452049 350829
rect 451813 350273 452049 350509
rect 467952 350593 468188 350829
rect 467952 350273 468188 350509
rect 473882 350593 474118 350829
rect 473882 350273 474118 350509
rect 479813 350593 480049 350829
rect 479813 350273 480049 350509
rect 495952 350593 496188 350829
rect 495952 350273 496188 350509
rect 501882 350593 502118 350829
rect 501882 350273 502118 350509
rect 507813 350593 508049 350829
rect 507813 350273 508049 350509
rect 523952 350593 524188 350829
rect 523952 350273 524188 350509
rect 529882 350593 530118 350829
rect 529882 350273 530118 350509
rect 535813 350593 536049 350829
rect 535813 350273 536049 350509
rect 551952 350593 552188 350829
rect 551952 350273 552188 350509
rect 557882 350593 558118 350829
rect 557882 350273 558118 350509
rect 563813 350593 564049 350829
rect 563813 350273 564049 350509
rect 573526 350593 573762 350829
rect 573846 350593 574082 350829
rect 573526 350273 573762 350509
rect 573846 350273 574082 350509
rect 22916 347218 23152 347454
rect 22916 346898 23152 347134
rect 28847 347218 29083 347454
rect 28847 346898 29083 347134
rect 50916 347218 51152 347454
rect 50916 346898 51152 347134
rect 56847 347218 57083 347454
rect 56847 346898 57083 347134
rect 78916 347218 79152 347454
rect 78916 346898 79152 347134
rect 84847 347218 85083 347454
rect 84847 346898 85083 347134
rect 106916 347218 107152 347454
rect 106916 346898 107152 347134
rect 112847 347218 113083 347454
rect 112847 346898 113083 347134
rect 134916 347218 135152 347454
rect 134916 346898 135152 347134
rect 140847 347218 141083 347454
rect 140847 346898 141083 347134
rect 162916 347218 163152 347454
rect 162916 346898 163152 347134
rect 168847 347218 169083 347454
rect 168847 346898 169083 347134
rect 190916 347218 191152 347454
rect 190916 346898 191152 347134
rect 196847 347218 197083 347454
rect 196847 346898 197083 347134
rect 218916 347218 219152 347454
rect 218916 346898 219152 347134
rect 224847 347218 225083 347454
rect 224847 346898 225083 347134
rect 246916 347218 247152 347454
rect 246916 346898 247152 347134
rect 252847 347218 253083 347454
rect 252847 346898 253083 347134
rect 274916 347218 275152 347454
rect 274916 346898 275152 347134
rect 280847 347218 281083 347454
rect 280847 346898 281083 347134
rect 302916 347218 303152 347454
rect 302916 346898 303152 347134
rect 308847 347218 309083 347454
rect 308847 346898 309083 347134
rect 330916 347218 331152 347454
rect 330916 346898 331152 347134
rect 336847 347218 337083 347454
rect 336847 346898 337083 347134
rect 358916 347218 359152 347454
rect 358916 346898 359152 347134
rect 364847 347218 365083 347454
rect 364847 346898 365083 347134
rect 386916 347218 387152 347454
rect 386916 346898 387152 347134
rect 392847 347218 393083 347454
rect 392847 346898 393083 347134
rect 414916 347218 415152 347454
rect 414916 346898 415152 347134
rect 420847 347218 421083 347454
rect 420847 346898 421083 347134
rect 442916 347218 443152 347454
rect 442916 346898 443152 347134
rect 448847 347218 449083 347454
rect 448847 346898 449083 347134
rect 470916 347218 471152 347454
rect 470916 346898 471152 347134
rect 476847 347218 477083 347454
rect 476847 346898 477083 347134
rect 498916 347218 499152 347454
rect 498916 346898 499152 347134
rect 504847 347218 505083 347454
rect 504847 346898 505083 347134
rect 526916 347218 527152 347454
rect 526916 346898 527152 347134
rect 532847 347218 533083 347454
rect 532847 346898 533083 347134
rect 554916 347218 555152 347454
rect 554916 346898 555152 347134
rect 560847 347218 561083 347454
rect 560847 346898 561083 347134
rect -1974 323593 -1738 323829
rect -1654 323593 -1418 323829
rect -1974 323273 -1738 323509
rect -1654 323273 -1418 323509
rect 19952 323593 20188 323829
rect 19952 323273 20188 323509
rect 25882 323593 26118 323829
rect 25882 323273 26118 323509
rect 31813 323593 32049 323829
rect 31813 323273 32049 323509
rect 47952 323593 48188 323829
rect 47952 323273 48188 323509
rect 53882 323593 54118 323829
rect 53882 323273 54118 323509
rect 59813 323593 60049 323829
rect 59813 323273 60049 323509
rect 75952 323593 76188 323829
rect 75952 323273 76188 323509
rect 81882 323593 82118 323829
rect 81882 323273 82118 323509
rect 87813 323593 88049 323829
rect 87813 323273 88049 323509
rect 103952 323593 104188 323829
rect 103952 323273 104188 323509
rect 109882 323593 110118 323829
rect 109882 323273 110118 323509
rect 115813 323593 116049 323829
rect 115813 323273 116049 323509
rect 131952 323593 132188 323829
rect 131952 323273 132188 323509
rect 137882 323593 138118 323829
rect 137882 323273 138118 323509
rect 143813 323593 144049 323829
rect 143813 323273 144049 323509
rect 159952 323593 160188 323829
rect 159952 323273 160188 323509
rect 165882 323593 166118 323829
rect 165882 323273 166118 323509
rect 171813 323593 172049 323829
rect 171813 323273 172049 323509
rect 187952 323593 188188 323829
rect 187952 323273 188188 323509
rect 193882 323593 194118 323829
rect 193882 323273 194118 323509
rect 199813 323593 200049 323829
rect 199813 323273 200049 323509
rect 215952 323593 216188 323829
rect 215952 323273 216188 323509
rect 221882 323593 222118 323829
rect 221882 323273 222118 323509
rect 227813 323593 228049 323829
rect 227813 323273 228049 323509
rect 243952 323593 244188 323829
rect 243952 323273 244188 323509
rect 249882 323593 250118 323829
rect 249882 323273 250118 323509
rect 255813 323593 256049 323829
rect 255813 323273 256049 323509
rect 271952 323593 272188 323829
rect 271952 323273 272188 323509
rect 277882 323593 278118 323829
rect 277882 323273 278118 323509
rect 283813 323593 284049 323829
rect 283813 323273 284049 323509
rect 299952 323593 300188 323829
rect 299952 323273 300188 323509
rect 305882 323593 306118 323829
rect 305882 323273 306118 323509
rect 311813 323593 312049 323829
rect 311813 323273 312049 323509
rect 327952 323593 328188 323829
rect 327952 323273 328188 323509
rect 333882 323593 334118 323829
rect 333882 323273 334118 323509
rect 339813 323593 340049 323829
rect 339813 323273 340049 323509
rect 355952 323593 356188 323829
rect 355952 323273 356188 323509
rect 361882 323593 362118 323829
rect 361882 323273 362118 323509
rect 367813 323593 368049 323829
rect 367813 323273 368049 323509
rect 383952 323593 384188 323829
rect 383952 323273 384188 323509
rect 389882 323593 390118 323829
rect 389882 323273 390118 323509
rect 395813 323593 396049 323829
rect 395813 323273 396049 323509
rect 411952 323593 412188 323829
rect 411952 323273 412188 323509
rect 417882 323593 418118 323829
rect 417882 323273 418118 323509
rect 423813 323593 424049 323829
rect 423813 323273 424049 323509
rect 439952 323593 440188 323829
rect 439952 323273 440188 323509
rect 445882 323593 446118 323829
rect 445882 323273 446118 323509
rect 451813 323593 452049 323829
rect 451813 323273 452049 323509
rect 467952 323593 468188 323829
rect 467952 323273 468188 323509
rect 473882 323593 474118 323829
rect 473882 323273 474118 323509
rect 479813 323593 480049 323829
rect 479813 323273 480049 323509
rect 495952 323593 496188 323829
rect 495952 323273 496188 323509
rect 501882 323593 502118 323829
rect 501882 323273 502118 323509
rect 507813 323593 508049 323829
rect 507813 323273 508049 323509
rect 523952 323593 524188 323829
rect 523952 323273 524188 323509
rect 529882 323593 530118 323829
rect 529882 323273 530118 323509
rect 535813 323593 536049 323829
rect 535813 323273 536049 323509
rect 551952 323593 552188 323829
rect 551952 323273 552188 323509
rect 557882 323593 558118 323829
rect 557882 323273 558118 323509
rect 563813 323593 564049 323829
rect 563813 323273 564049 323509
rect 573526 323593 573762 323829
rect 573846 323593 574082 323829
rect 573526 323273 573762 323509
rect 573846 323273 574082 323509
rect 22916 320218 23152 320454
rect 22916 319898 23152 320134
rect 28847 320218 29083 320454
rect 28847 319898 29083 320134
rect 50916 320218 51152 320454
rect 50916 319898 51152 320134
rect 56847 320218 57083 320454
rect 56847 319898 57083 320134
rect 78916 320218 79152 320454
rect 78916 319898 79152 320134
rect 84847 320218 85083 320454
rect 84847 319898 85083 320134
rect 106916 320218 107152 320454
rect 106916 319898 107152 320134
rect 112847 320218 113083 320454
rect 112847 319898 113083 320134
rect 134916 320218 135152 320454
rect 134916 319898 135152 320134
rect 140847 320218 141083 320454
rect 140847 319898 141083 320134
rect 162916 320218 163152 320454
rect 162916 319898 163152 320134
rect 168847 320218 169083 320454
rect 168847 319898 169083 320134
rect 190916 320218 191152 320454
rect 190916 319898 191152 320134
rect 196847 320218 197083 320454
rect 196847 319898 197083 320134
rect 218916 320218 219152 320454
rect 218916 319898 219152 320134
rect 224847 320218 225083 320454
rect 224847 319898 225083 320134
rect 246916 320218 247152 320454
rect 246916 319898 247152 320134
rect 252847 320218 253083 320454
rect 252847 319898 253083 320134
rect 274916 320218 275152 320454
rect 274916 319898 275152 320134
rect 280847 320218 281083 320454
rect 280847 319898 281083 320134
rect 302916 320218 303152 320454
rect 302916 319898 303152 320134
rect 308847 320218 309083 320454
rect 308847 319898 309083 320134
rect 330916 320218 331152 320454
rect 330916 319898 331152 320134
rect 336847 320218 337083 320454
rect 336847 319898 337083 320134
rect 358916 320218 359152 320454
rect 358916 319898 359152 320134
rect 364847 320218 365083 320454
rect 364847 319898 365083 320134
rect 386916 320218 387152 320454
rect 386916 319898 387152 320134
rect 392847 320218 393083 320454
rect 392847 319898 393083 320134
rect 414916 320218 415152 320454
rect 414916 319898 415152 320134
rect 420847 320218 421083 320454
rect 420847 319898 421083 320134
rect 442916 320218 443152 320454
rect 442916 319898 443152 320134
rect 448847 320218 449083 320454
rect 448847 319898 449083 320134
rect 470916 320218 471152 320454
rect 470916 319898 471152 320134
rect 476847 320218 477083 320454
rect 476847 319898 477083 320134
rect 498916 320218 499152 320454
rect 498916 319898 499152 320134
rect 504847 320218 505083 320454
rect 504847 319898 505083 320134
rect 526916 320218 527152 320454
rect 526916 319898 527152 320134
rect 532847 320218 533083 320454
rect 532847 319898 533083 320134
rect 554916 320218 555152 320454
rect 554916 319898 555152 320134
rect 560847 320218 561083 320454
rect 560847 319898 561083 320134
rect -1974 296593 -1738 296829
rect -1654 296593 -1418 296829
rect -1974 296273 -1738 296509
rect -1654 296273 -1418 296509
rect 19952 296593 20188 296829
rect 19952 296273 20188 296509
rect 25882 296593 26118 296829
rect 25882 296273 26118 296509
rect 31813 296593 32049 296829
rect 31813 296273 32049 296509
rect 47952 296593 48188 296829
rect 47952 296273 48188 296509
rect 53882 296593 54118 296829
rect 53882 296273 54118 296509
rect 59813 296593 60049 296829
rect 59813 296273 60049 296509
rect 75952 296593 76188 296829
rect 75952 296273 76188 296509
rect 81882 296593 82118 296829
rect 81882 296273 82118 296509
rect 87813 296593 88049 296829
rect 87813 296273 88049 296509
rect 103952 296593 104188 296829
rect 103952 296273 104188 296509
rect 109882 296593 110118 296829
rect 109882 296273 110118 296509
rect 115813 296593 116049 296829
rect 115813 296273 116049 296509
rect 131952 296593 132188 296829
rect 131952 296273 132188 296509
rect 137882 296593 138118 296829
rect 137882 296273 138118 296509
rect 143813 296593 144049 296829
rect 143813 296273 144049 296509
rect 159952 296593 160188 296829
rect 159952 296273 160188 296509
rect 165882 296593 166118 296829
rect 165882 296273 166118 296509
rect 171813 296593 172049 296829
rect 171813 296273 172049 296509
rect 187952 296593 188188 296829
rect 187952 296273 188188 296509
rect 193882 296593 194118 296829
rect 193882 296273 194118 296509
rect 199813 296593 200049 296829
rect 199813 296273 200049 296509
rect 215952 296593 216188 296829
rect 215952 296273 216188 296509
rect 221882 296593 222118 296829
rect 221882 296273 222118 296509
rect 227813 296593 228049 296829
rect 227813 296273 228049 296509
rect 243952 296593 244188 296829
rect 243952 296273 244188 296509
rect 249882 296593 250118 296829
rect 249882 296273 250118 296509
rect 255813 296593 256049 296829
rect 255813 296273 256049 296509
rect 271952 296593 272188 296829
rect 271952 296273 272188 296509
rect 277882 296593 278118 296829
rect 277882 296273 278118 296509
rect 283813 296593 284049 296829
rect 283813 296273 284049 296509
rect 299952 296593 300188 296829
rect 299952 296273 300188 296509
rect 305882 296593 306118 296829
rect 305882 296273 306118 296509
rect 311813 296593 312049 296829
rect 311813 296273 312049 296509
rect 327952 296593 328188 296829
rect 327952 296273 328188 296509
rect 333882 296593 334118 296829
rect 333882 296273 334118 296509
rect 339813 296593 340049 296829
rect 339813 296273 340049 296509
rect 355952 296593 356188 296829
rect 355952 296273 356188 296509
rect 361882 296593 362118 296829
rect 361882 296273 362118 296509
rect 367813 296593 368049 296829
rect 367813 296273 368049 296509
rect 383952 296593 384188 296829
rect 383952 296273 384188 296509
rect 389882 296593 390118 296829
rect 389882 296273 390118 296509
rect 395813 296593 396049 296829
rect 395813 296273 396049 296509
rect 411952 296593 412188 296829
rect 411952 296273 412188 296509
rect 417882 296593 418118 296829
rect 417882 296273 418118 296509
rect 423813 296593 424049 296829
rect 423813 296273 424049 296509
rect 439952 296593 440188 296829
rect 439952 296273 440188 296509
rect 445882 296593 446118 296829
rect 445882 296273 446118 296509
rect 451813 296593 452049 296829
rect 451813 296273 452049 296509
rect 467952 296593 468188 296829
rect 467952 296273 468188 296509
rect 473882 296593 474118 296829
rect 473882 296273 474118 296509
rect 479813 296593 480049 296829
rect 479813 296273 480049 296509
rect 495952 296593 496188 296829
rect 495952 296273 496188 296509
rect 501882 296593 502118 296829
rect 501882 296273 502118 296509
rect 507813 296593 508049 296829
rect 507813 296273 508049 296509
rect 523952 296593 524188 296829
rect 523952 296273 524188 296509
rect 529882 296593 530118 296829
rect 529882 296273 530118 296509
rect 535813 296593 536049 296829
rect 535813 296273 536049 296509
rect 551952 296593 552188 296829
rect 551952 296273 552188 296509
rect 557882 296593 558118 296829
rect 557882 296273 558118 296509
rect 563813 296593 564049 296829
rect 563813 296273 564049 296509
rect 573526 296593 573762 296829
rect 573846 296593 574082 296829
rect 573526 296273 573762 296509
rect 573846 296273 574082 296509
rect 22916 293218 23152 293454
rect 22916 292898 23152 293134
rect 28847 293218 29083 293454
rect 28847 292898 29083 293134
rect 50916 293218 51152 293454
rect 50916 292898 51152 293134
rect 56847 293218 57083 293454
rect 56847 292898 57083 293134
rect 78916 293218 79152 293454
rect 78916 292898 79152 293134
rect 84847 293218 85083 293454
rect 84847 292898 85083 293134
rect 106916 293218 107152 293454
rect 106916 292898 107152 293134
rect 112847 293218 113083 293454
rect 112847 292898 113083 293134
rect 134916 293218 135152 293454
rect 134916 292898 135152 293134
rect 140847 293218 141083 293454
rect 140847 292898 141083 293134
rect 162916 293218 163152 293454
rect 162916 292898 163152 293134
rect 168847 293218 169083 293454
rect 168847 292898 169083 293134
rect 190916 293218 191152 293454
rect 190916 292898 191152 293134
rect 196847 293218 197083 293454
rect 196847 292898 197083 293134
rect 218916 293218 219152 293454
rect 218916 292898 219152 293134
rect 224847 293218 225083 293454
rect 224847 292898 225083 293134
rect 246916 293218 247152 293454
rect 246916 292898 247152 293134
rect 252847 293218 253083 293454
rect 252847 292898 253083 293134
rect 274916 293218 275152 293454
rect 274916 292898 275152 293134
rect 280847 293218 281083 293454
rect 280847 292898 281083 293134
rect 302916 293218 303152 293454
rect 302916 292898 303152 293134
rect 308847 293218 309083 293454
rect 308847 292898 309083 293134
rect 330916 293218 331152 293454
rect 330916 292898 331152 293134
rect 336847 293218 337083 293454
rect 336847 292898 337083 293134
rect 358916 293218 359152 293454
rect 358916 292898 359152 293134
rect 364847 293218 365083 293454
rect 364847 292898 365083 293134
rect 386916 293218 387152 293454
rect 386916 292898 387152 293134
rect 392847 293218 393083 293454
rect 392847 292898 393083 293134
rect 414916 293218 415152 293454
rect 414916 292898 415152 293134
rect 420847 293218 421083 293454
rect 420847 292898 421083 293134
rect 442916 293218 443152 293454
rect 442916 292898 443152 293134
rect 448847 293218 449083 293454
rect 448847 292898 449083 293134
rect 470916 293218 471152 293454
rect 470916 292898 471152 293134
rect 476847 293218 477083 293454
rect 476847 292898 477083 293134
rect 498916 293218 499152 293454
rect 498916 292898 499152 293134
rect 504847 293218 505083 293454
rect 504847 292898 505083 293134
rect 526916 293218 527152 293454
rect 526916 292898 527152 293134
rect 532847 293218 533083 293454
rect 532847 292898 533083 293134
rect 554916 293218 555152 293454
rect 554916 292898 555152 293134
rect 560847 293218 561083 293454
rect 560847 292898 561083 293134
rect -1974 269593 -1738 269829
rect -1654 269593 -1418 269829
rect -1974 269273 -1738 269509
rect -1654 269273 -1418 269509
rect 19952 269593 20188 269829
rect 19952 269273 20188 269509
rect 25882 269593 26118 269829
rect 25882 269273 26118 269509
rect 31813 269593 32049 269829
rect 31813 269273 32049 269509
rect 47952 269593 48188 269829
rect 47952 269273 48188 269509
rect 53882 269593 54118 269829
rect 53882 269273 54118 269509
rect 59813 269593 60049 269829
rect 59813 269273 60049 269509
rect 75952 269593 76188 269829
rect 75952 269273 76188 269509
rect 81882 269593 82118 269829
rect 81882 269273 82118 269509
rect 87813 269593 88049 269829
rect 87813 269273 88049 269509
rect 103952 269593 104188 269829
rect 103952 269273 104188 269509
rect 109882 269593 110118 269829
rect 109882 269273 110118 269509
rect 115813 269593 116049 269829
rect 115813 269273 116049 269509
rect 131952 269593 132188 269829
rect 131952 269273 132188 269509
rect 137882 269593 138118 269829
rect 137882 269273 138118 269509
rect 143813 269593 144049 269829
rect 143813 269273 144049 269509
rect 159952 269593 160188 269829
rect 159952 269273 160188 269509
rect 165882 269593 166118 269829
rect 165882 269273 166118 269509
rect 171813 269593 172049 269829
rect 171813 269273 172049 269509
rect 187952 269593 188188 269829
rect 187952 269273 188188 269509
rect 193882 269593 194118 269829
rect 193882 269273 194118 269509
rect 199813 269593 200049 269829
rect 199813 269273 200049 269509
rect 215952 269593 216188 269829
rect 215952 269273 216188 269509
rect 221882 269593 222118 269829
rect 221882 269273 222118 269509
rect 227813 269593 228049 269829
rect 227813 269273 228049 269509
rect 243952 269593 244188 269829
rect 243952 269273 244188 269509
rect 249882 269593 250118 269829
rect 249882 269273 250118 269509
rect 255813 269593 256049 269829
rect 255813 269273 256049 269509
rect 271952 269593 272188 269829
rect 271952 269273 272188 269509
rect 277882 269593 278118 269829
rect 277882 269273 278118 269509
rect 283813 269593 284049 269829
rect 283813 269273 284049 269509
rect 299952 269593 300188 269829
rect 299952 269273 300188 269509
rect 305882 269593 306118 269829
rect 305882 269273 306118 269509
rect 311813 269593 312049 269829
rect 311813 269273 312049 269509
rect 327952 269593 328188 269829
rect 327952 269273 328188 269509
rect 333882 269593 334118 269829
rect 333882 269273 334118 269509
rect 339813 269593 340049 269829
rect 339813 269273 340049 269509
rect 355952 269593 356188 269829
rect 355952 269273 356188 269509
rect 361882 269593 362118 269829
rect 361882 269273 362118 269509
rect 367813 269593 368049 269829
rect 367813 269273 368049 269509
rect 383952 269593 384188 269829
rect 383952 269273 384188 269509
rect 389882 269593 390118 269829
rect 389882 269273 390118 269509
rect 395813 269593 396049 269829
rect 395813 269273 396049 269509
rect 411952 269593 412188 269829
rect 411952 269273 412188 269509
rect 417882 269593 418118 269829
rect 417882 269273 418118 269509
rect 423813 269593 424049 269829
rect 423813 269273 424049 269509
rect 439952 269593 440188 269829
rect 439952 269273 440188 269509
rect 445882 269593 446118 269829
rect 445882 269273 446118 269509
rect 451813 269593 452049 269829
rect 451813 269273 452049 269509
rect 467952 269593 468188 269829
rect 467952 269273 468188 269509
rect 473882 269593 474118 269829
rect 473882 269273 474118 269509
rect 479813 269593 480049 269829
rect 479813 269273 480049 269509
rect 495952 269593 496188 269829
rect 495952 269273 496188 269509
rect 501882 269593 502118 269829
rect 501882 269273 502118 269509
rect 507813 269593 508049 269829
rect 507813 269273 508049 269509
rect 523952 269593 524188 269829
rect 523952 269273 524188 269509
rect 529882 269593 530118 269829
rect 529882 269273 530118 269509
rect 535813 269593 536049 269829
rect 535813 269273 536049 269509
rect 551952 269593 552188 269829
rect 551952 269273 552188 269509
rect 557882 269593 558118 269829
rect 557882 269273 558118 269509
rect 563813 269593 564049 269829
rect 563813 269273 564049 269509
rect 573526 269593 573762 269829
rect 573846 269593 574082 269829
rect 573526 269273 573762 269509
rect 573846 269273 574082 269509
rect 22916 266218 23152 266454
rect 22916 265898 23152 266134
rect 28847 266218 29083 266454
rect 28847 265898 29083 266134
rect 50916 266218 51152 266454
rect 50916 265898 51152 266134
rect 56847 266218 57083 266454
rect 56847 265898 57083 266134
rect 78916 266218 79152 266454
rect 78916 265898 79152 266134
rect 84847 266218 85083 266454
rect 84847 265898 85083 266134
rect 106916 266218 107152 266454
rect 106916 265898 107152 266134
rect 112847 266218 113083 266454
rect 112847 265898 113083 266134
rect 134916 266218 135152 266454
rect 134916 265898 135152 266134
rect 140847 266218 141083 266454
rect 140847 265898 141083 266134
rect 162916 266218 163152 266454
rect 162916 265898 163152 266134
rect 168847 266218 169083 266454
rect 168847 265898 169083 266134
rect 190916 266218 191152 266454
rect 190916 265898 191152 266134
rect 196847 266218 197083 266454
rect 196847 265898 197083 266134
rect 218916 266218 219152 266454
rect 218916 265898 219152 266134
rect 224847 266218 225083 266454
rect 224847 265898 225083 266134
rect 246916 266218 247152 266454
rect 246916 265898 247152 266134
rect 252847 266218 253083 266454
rect 252847 265898 253083 266134
rect 274916 266218 275152 266454
rect 274916 265898 275152 266134
rect 280847 266218 281083 266454
rect 280847 265898 281083 266134
rect 302916 266218 303152 266454
rect 302916 265898 303152 266134
rect 308847 266218 309083 266454
rect 308847 265898 309083 266134
rect 330916 266218 331152 266454
rect 330916 265898 331152 266134
rect 336847 266218 337083 266454
rect 336847 265898 337083 266134
rect 358916 266218 359152 266454
rect 358916 265898 359152 266134
rect 364847 266218 365083 266454
rect 364847 265898 365083 266134
rect 386916 266218 387152 266454
rect 386916 265898 387152 266134
rect 392847 266218 393083 266454
rect 392847 265898 393083 266134
rect 414916 266218 415152 266454
rect 414916 265898 415152 266134
rect 420847 266218 421083 266454
rect 420847 265898 421083 266134
rect 442916 266218 443152 266454
rect 442916 265898 443152 266134
rect 448847 266218 449083 266454
rect 448847 265898 449083 266134
rect 470916 266218 471152 266454
rect 470916 265898 471152 266134
rect 476847 266218 477083 266454
rect 476847 265898 477083 266134
rect 498916 266218 499152 266454
rect 498916 265898 499152 266134
rect 504847 266218 505083 266454
rect 504847 265898 505083 266134
rect 526916 266218 527152 266454
rect 526916 265898 527152 266134
rect 532847 266218 533083 266454
rect 532847 265898 533083 266134
rect 554916 266218 555152 266454
rect 554916 265898 555152 266134
rect 560847 266218 561083 266454
rect 560847 265898 561083 266134
rect -1974 242593 -1738 242829
rect -1654 242593 -1418 242829
rect -1974 242273 -1738 242509
rect -1654 242273 -1418 242509
rect 19952 242593 20188 242829
rect 19952 242273 20188 242509
rect 25882 242593 26118 242829
rect 25882 242273 26118 242509
rect 31813 242593 32049 242829
rect 31813 242273 32049 242509
rect 47952 242593 48188 242829
rect 47952 242273 48188 242509
rect 53882 242593 54118 242829
rect 53882 242273 54118 242509
rect 59813 242593 60049 242829
rect 59813 242273 60049 242509
rect 75952 242593 76188 242829
rect 75952 242273 76188 242509
rect 81882 242593 82118 242829
rect 81882 242273 82118 242509
rect 87813 242593 88049 242829
rect 87813 242273 88049 242509
rect 103952 242593 104188 242829
rect 103952 242273 104188 242509
rect 109882 242593 110118 242829
rect 109882 242273 110118 242509
rect 115813 242593 116049 242829
rect 115813 242273 116049 242509
rect 131952 242593 132188 242829
rect 131952 242273 132188 242509
rect 137882 242593 138118 242829
rect 137882 242273 138118 242509
rect 143813 242593 144049 242829
rect 143813 242273 144049 242509
rect 159952 242593 160188 242829
rect 159952 242273 160188 242509
rect 165882 242593 166118 242829
rect 165882 242273 166118 242509
rect 171813 242593 172049 242829
rect 171813 242273 172049 242509
rect 187952 242593 188188 242829
rect 187952 242273 188188 242509
rect 193882 242593 194118 242829
rect 193882 242273 194118 242509
rect 199813 242593 200049 242829
rect 199813 242273 200049 242509
rect 215952 242593 216188 242829
rect 215952 242273 216188 242509
rect 221882 242593 222118 242829
rect 221882 242273 222118 242509
rect 227813 242593 228049 242829
rect 227813 242273 228049 242509
rect 243952 242593 244188 242829
rect 243952 242273 244188 242509
rect 249882 242593 250118 242829
rect 249882 242273 250118 242509
rect 255813 242593 256049 242829
rect 255813 242273 256049 242509
rect 271952 242593 272188 242829
rect 271952 242273 272188 242509
rect 277882 242593 278118 242829
rect 277882 242273 278118 242509
rect 283813 242593 284049 242829
rect 283813 242273 284049 242509
rect 299952 242593 300188 242829
rect 299952 242273 300188 242509
rect 305882 242593 306118 242829
rect 305882 242273 306118 242509
rect 311813 242593 312049 242829
rect 311813 242273 312049 242509
rect 327952 242593 328188 242829
rect 327952 242273 328188 242509
rect 333882 242593 334118 242829
rect 333882 242273 334118 242509
rect 339813 242593 340049 242829
rect 339813 242273 340049 242509
rect 355952 242593 356188 242829
rect 355952 242273 356188 242509
rect 361882 242593 362118 242829
rect 361882 242273 362118 242509
rect 367813 242593 368049 242829
rect 367813 242273 368049 242509
rect 383952 242593 384188 242829
rect 383952 242273 384188 242509
rect 389882 242593 390118 242829
rect 389882 242273 390118 242509
rect 395813 242593 396049 242829
rect 395813 242273 396049 242509
rect 411952 242593 412188 242829
rect 411952 242273 412188 242509
rect 417882 242593 418118 242829
rect 417882 242273 418118 242509
rect 423813 242593 424049 242829
rect 423813 242273 424049 242509
rect 439952 242593 440188 242829
rect 439952 242273 440188 242509
rect 445882 242593 446118 242829
rect 445882 242273 446118 242509
rect 451813 242593 452049 242829
rect 451813 242273 452049 242509
rect 467952 242593 468188 242829
rect 467952 242273 468188 242509
rect 473882 242593 474118 242829
rect 473882 242273 474118 242509
rect 479813 242593 480049 242829
rect 479813 242273 480049 242509
rect 495952 242593 496188 242829
rect 495952 242273 496188 242509
rect 501882 242593 502118 242829
rect 501882 242273 502118 242509
rect 507813 242593 508049 242829
rect 507813 242273 508049 242509
rect 523952 242593 524188 242829
rect 523952 242273 524188 242509
rect 529882 242593 530118 242829
rect 529882 242273 530118 242509
rect 535813 242593 536049 242829
rect 535813 242273 536049 242509
rect 551952 242593 552188 242829
rect 551952 242273 552188 242509
rect 557882 242593 558118 242829
rect 557882 242273 558118 242509
rect 563813 242593 564049 242829
rect 563813 242273 564049 242509
rect 573526 242593 573762 242829
rect 573846 242593 574082 242829
rect 573526 242273 573762 242509
rect 573846 242273 574082 242509
rect 22916 239218 23152 239454
rect 22916 238898 23152 239134
rect 28847 239218 29083 239454
rect 28847 238898 29083 239134
rect 50916 239218 51152 239454
rect 50916 238898 51152 239134
rect 56847 239218 57083 239454
rect 56847 238898 57083 239134
rect 78916 239218 79152 239454
rect 78916 238898 79152 239134
rect 84847 239218 85083 239454
rect 84847 238898 85083 239134
rect 106916 239218 107152 239454
rect 106916 238898 107152 239134
rect 112847 239218 113083 239454
rect 112847 238898 113083 239134
rect 134916 239218 135152 239454
rect 134916 238898 135152 239134
rect 140847 239218 141083 239454
rect 140847 238898 141083 239134
rect 162916 239218 163152 239454
rect 162916 238898 163152 239134
rect 168847 239218 169083 239454
rect 168847 238898 169083 239134
rect 190916 239218 191152 239454
rect 190916 238898 191152 239134
rect 196847 239218 197083 239454
rect 196847 238898 197083 239134
rect 218916 239218 219152 239454
rect 218916 238898 219152 239134
rect 224847 239218 225083 239454
rect 224847 238898 225083 239134
rect 246916 239218 247152 239454
rect 246916 238898 247152 239134
rect 252847 239218 253083 239454
rect 252847 238898 253083 239134
rect 274916 239218 275152 239454
rect 274916 238898 275152 239134
rect 280847 239218 281083 239454
rect 280847 238898 281083 239134
rect 302916 239218 303152 239454
rect 302916 238898 303152 239134
rect 308847 239218 309083 239454
rect 308847 238898 309083 239134
rect 330916 239218 331152 239454
rect 330916 238898 331152 239134
rect 336847 239218 337083 239454
rect 336847 238898 337083 239134
rect 358916 239218 359152 239454
rect 358916 238898 359152 239134
rect 364847 239218 365083 239454
rect 364847 238898 365083 239134
rect 386916 239218 387152 239454
rect 386916 238898 387152 239134
rect 392847 239218 393083 239454
rect 392847 238898 393083 239134
rect 414916 239218 415152 239454
rect 414916 238898 415152 239134
rect 420847 239218 421083 239454
rect 420847 238898 421083 239134
rect 442916 239218 443152 239454
rect 442916 238898 443152 239134
rect 448847 239218 449083 239454
rect 448847 238898 449083 239134
rect 470916 239218 471152 239454
rect 470916 238898 471152 239134
rect 476847 239218 477083 239454
rect 476847 238898 477083 239134
rect 498916 239218 499152 239454
rect 498916 238898 499152 239134
rect 504847 239218 505083 239454
rect 504847 238898 505083 239134
rect 526916 239218 527152 239454
rect 526916 238898 527152 239134
rect 532847 239218 533083 239454
rect 532847 238898 533083 239134
rect 554916 239218 555152 239454
rect 554916 238898 555152 239134
rect 560847 239218 561083 239454
rect 560847 238898 561083 239134
rect -1974 215593 -1738 215829
rect -1654 215593 -1418 215829
rect -1974 215273 -1738 215509
rect -1654 215273 -1418 215509
rect 19952 215593 20188 215829
rect 19952 215273 20188 215509
rect 25882 215593 26118 215829
rect 25882 215273 26118 215509
rect 31813 215593 32049 215829
rect 31813 215273 32049 215509
rect 47952 215593 48188 215829
rect 47952 215273 48188 215509
rect 53882 215593 54118 215829
rect 53882 215273 54118 215509
rect 59813 215593 60049 215829
rect 59813 215273 60049 215509
rect 75952 215593 76188 215829
rect 75952 215273 76188 215509
rect 81882 215593 82118 215829
rect 81882 215273 82118 215509
rect 87813 215593 88049 215829
rect 87813 215273 88049 215509
rect 103952 215593 104188 215829
rect 103952 215273 104188 215509
rect 109882 215593 110118 215829
rect 109882 215273 110118 215509
rect 115813 215593 116049 215829
rect 115813 215273 116049 215509
rect 131952 215593 132188 215829
rect 131952 215273 132188 215509
rect 137882 215593 138118 215829
rect 137882 215273 138118 215509
rect 143813 215593 144049 215829
rect 143813 215273 144049 215509
rect 159952 215593 160188 215829
rect 159952 215273 160188 215509
rect 165882 215593 166118 215829
rect 165882 215273 166118 215509
rect 171813 215593 172049 215829
rect 171813 215273 172049 215509
rect 187952 215593 188188 215829
rect 187952 215273 188188 215509
rect 193882 215593 194118 215829
rect 193882 215273 194118 215509
rect 199813 215593 200049 215829
rect 199813 215273 200049 215509
rect 215952 215593 216188 215829
rect 215952 215273 216188 215509
rect 221882 215593 222118 215829
rect 221882 215273 222118 215509
rect 227813 215593 228049 215829
rect 227813 215273 228049 215509
rect 243952 215593 244188 215829
rect 243952 215273 244188 215509
rect 249882 215593 250118 215829
rect 249882 215273 250118 215509
rect 255813 215593 256049 215829
rect 255813 215273 256049 215509
rect 271952 215593 272188 215829
rect 271952 215273 272188 215509
rect 277882 215593 278118 215829
rect 277882 215273 278118 215509
rect 283813 215593 284049 215829
rect 283813 215273 284049 215509
rect 299952 215593 300188 215829
rect 299952 215273 300188 215509
rect 305882 215593 306118 215829
rect 305882 215273 306118 215509
rect 311813 215593 312049 215829
rect 311813 215273 312049 215509
rect 327952 215593 328188 215829
rect 327952 215273 328188 215509
rect 333882 215593 334118 215829
rect 333882 215273 334118 215509
rect 339813 215593 340049 215829
rect 339813 215273 340049 215509
rect 355952 215593 356188 215829
rect 355952 215273 356188 215509
rect 361882 215593 362118 215829
rect 361882 215273 362118 215509
rect 367813 215593 368049 215829
rect 367813 215273 368049 215509
rect 383952 215593 384188 215829
rect 383952 215273 384188 215509
rect 389882 215593 390118 215829
rect 389882 215273 390118 215509
rect 395813 215593 396049 215829
rect 395813 215273 396049 215509
rect 411952 215593 412188 215829
rect 411952 215273 412188 215509
rect 417882 215593 418118 215829
rect 417882 215273 418118 215509
rect 423813 215593 424049 215829
rect 423813 215273 424049 215509
rect 439952 215593 440188 215829
rect 439952 215273 440188 215509
rect 445882 215593 446118 215829
rect 445882 215273 446118 215509
rect 451813 215593 452049 215829
rect 451813 215273 452049 215509
rect 467952 215593 468188 215829
rect 467952 215273 468188 215509
rect 473882 215593 474118 215829
rect 473882 215273 474118 215509
rect 479813 215593 480049 215829
rect 479813 215273 480049 215509
rect 495952 215593 496188 215829
rect 495952 215273 496188 215509
rect 501882 215593 502118 215829
rect 501882 215273 502118 215509
rect 507813 215593 508049 215829
rect 507813 215273 508049 215509
rect 523952 215593 524188 215829
rect 523952 215273 524188 215509
rect 529882 215593 530118 215829
rect 529882 215273 530118 215509
rect 535813 215593 536049 215829
rect 535813 215273 536049 215509
rect 551952 215593 552188 215829
rect 551952 215273 552188 215509
rect 557882 215593 558118 215829
rect 557882 215273 558118 215509
rect 563813 215593 564049 215829
rect 563813 215273 564049 215509
rect 573526 215593 573762 215829
rect 573846 215593 574082 215829
rect 573526 215273 573762 215509
rect 573846 215273 574082 215509
rect 22916 212218 23152 212454
rect 22916 211898 23152 212134
rect 28847 212218 29083 212454
rect 28847 211898 29083 212134
rect 50916 212218 51152 212454
rect 50916 211898 51152 212134
rect 56847 212218 57083 212454
rect 56847 211898 57083 212134
rect 78916 212218 79152 212454
rect 78916 211898 79152 212134
rect 84847 212218 85083 212454
rect 84847 211898 85083 212134
rect 106916 212218 107152 212454
rect 106916 211898 107152 212134
rect 112847 212218 113083 212454
rect 112847 211898 113083 212134
rect 134916 212218 135152 212454
rect 134916 211898 135152 212134
rect 140847 212218 141083 212454
rect 140847 211898 141083 212134
rect 162916 212218 163152 212454
rect 162916 211898 163152 212134
rect 168847 212218 169083 212454
rect 168847 211898 169083 212134
rect 190916 212218 191152 212454
rect 190916 211898 191152 212134
rect 196847 212218 197083 212454
rect 196847 211898 197083 212134
rect 218916 212218 219152 212454
rect 218916 211898 219152 212134
rect 224847 212218 225083 212454
rect 224847 211898 225083 212134
rect 246916 212218 247152 212454
rect 246916 211898 247152 212134
rect 252847 212218 253083 212454
rect 252847 211898 253083 212134
rect 274916 212218 275152 212454
rect 274916 211898 275152 212134
rect 280847 212218 281083 212454
rect 280847 211898 281083 212134
rect 302916 212218 303152 212454
rect 302916 211898 303152 212134
rect 308847 212218 309083 212454
rect 308847 211898 309083 212134
rect 330916 212218 331152 212454
rect 330916 211898 331152 212134
rect 336847 212218 337083 212454
rect 336847 211898 337083 212134
rect 358916 212218 359152 212454
rect 358916 211898 359152 212134
rect 364847 212218 365083 212454
rect 364847 211898 365083 212134
rect 386916 212218 387152 212454
rect 386916 211898 387152 212134
rect 392847 212218 393083 212454
rect 392847 211898 393083 212134
rect 414916 212218 415152 212454
rect 414916 211898 415152 212134
rect 420847 212218 421083 212454
rect 420847 211898 421083 212134
rect 442916 212218 443152 212454
rect 442916 211898 443152 212134
rect 448847 212218 449083 212454
rect 448847 211898 449083 212134
rect 470916 212218 471152 212454
rect 470916 211898 471152 212134
rect 476847 212218 477083 212454
rect 476847 211898 477083 212134
rect 498916 212218 499152 212454
rect 498916 211898 499152 212134
rect 504847 212218 505083 212454
rect 504847 211898 505083 212134
rect 526916 212218 527152 212454
rect 526916 211898 527152 212134
rect 532847 212218 533083 212454
rect 532847 211898 533083 212134
rect 554916 212218 555152 212454
rect 554916 211898 555152 212134
rect 560847 212218 561083 212454
rect 560847 211898 561083 212134
rect -1974 188593 -1738 188829
rect -1654 188593 -1418 188829
rect -1974 188273 -1738 188509
rect -1654 188273 -1418 188509
rect 19952 188593 20188 188829
rect 19952 188273 20188 188509
rect 25882 188593 26118 188829
rect 25882 188273 26118 188509
rect 31813 188593 32049 188829
rect 31813 188273 32049 188509
rect 47952 188593 48188 188829
rect 47952 188273 48188 188509
rect 53882 188593 54118 188829
rect 53882 188273 54118 188509
rect 59813 188593 60049 188829
rect 59813 188273 60049 188509
rect 75952 188593 76188 188829
rect 75952 188273 76188 188509
rect 81882 188593 82118 188829
rect 81882 188273 82118 188509
rect 87813 188593 88049 188829
rect 87813 188273 88049 188509
rect 103952 188593 104188 188829
rect 103952 188273 104188 188509
rect 109882 188593 110118 188829
rect 109882 188273 110118 188509
rect 115813 188593 116049 188829
rect 115813 188273 116049 188509
rect 131952 188593 132188 188829
rect 131952 188273 132188 188509
rect 137882 188593 138118 188829
rect 137882 188273 138118 188509
rect 143813 188593 144049 188829
rect 143813 188273 144049 188509
rect 159952 188593 160188 188829
rect 159952 188273 160188 188509
rect 165882 188593 166118 188829
rect 165882 188273 166118 188509
rect 171813 188593 172049 188829
rect 171813 188273 172049 188509
rect 187952 188593 188188 188829
rect 187952 188273 188188 188509
rect 193882 188593 194118 188829
rect 193882 188273 194118 188509
rect 199813 188593 200049 188829
rect 199813 188273 200049 188509
rect 215952 188593 216188 188829
rect 215952 188273 216188 188509
rect 221882 188593 222118 188829
rect 221882 188273 222118 188509
rect 227813 188593 228049 188829
rect 227813 188273 228049 188509
rect 243952 188593 244188 188829
rect 243952 188273 244188 188509
rect 249882 188593 250118 188829
rect 249882 188273 250118 188509
rect 255813 188593 256049 188829
rect 255813 188273 256049 188509
rect 271952 188593 272188 188829
rect 271952 188273 272188 188509
rect 277882 188593 278118 188829
rect 277882 188273 278118 188509
rect 283813 188593 284049 188829
rect 283813 188273 284049 188509
rect 299952 188593 300188 188829
rect 299952 188273 300188 188509
rect 305882 188593 306118 188829
rect 305882 188273 306118 188509
rect 311813 188593 312049 188829
rect 311813 188273 312049 188509
rect 327952 188593 328188 188829
rect 327952 188273 328188 188509
rect 333882 188593 334118 188829
rect 333882 188273 334118 188509
rect 339813 188593 340049 188829
rect 339813 188273 340049 188509
rect 355952 188593 356188 188829
rect 355952 188273 356188 188509
rect 361882 188593 362118 188829
rect 361882 188273 362118 188509
rect 367813 188593 368049 188829
rect 367813 188273 368049 188509
rect 383952 188593 384188 188829
rect 383952 188273 384188 188509
rect 389882 188593 390118 188829
rect 389882 188273 390118 188509
rect 395813 188593 396049 188829
rect 395813 188273 396049 188509
rect 411952 188593 412188 188829
rect 411952 188273 412188 188509
rect 417882 188593 418118 188829
rect 417882 188273 418118 188509
rect 423813 188593 424049 188829
rect 423813 188273 424049 188509
rect 439952 188593 440188 188829
rect 439952 188273 440188 188509
rect 445882 188593 446118 188829
rect 445882 188273 446118 188509
rect 451813 188593 452049 188829
rect 451813 188273 452049 188509
rect 467952 188593 468188 188829
rect 467952 188273 468188 188509
rect 473882 188593 474118 188829
rect 473882 188273 474118 188509
rect 479813 188593 480049 188829
rect 479813 188273 480049 188509
rect 495952 188593 496188 188829
rect 495952 188273 496188 188509
rect 501882 188593 502118 188829
rect 501882 188273 502118 188509
rect 507813 188593 508049 188829
rect 507813 188273 508049 188509
rect 523952 188593 524188 188829
rect 523952 188273 524188 188509
rect 529882 188593 530118 188829
rect 529882 188273 530118 188509
rect 535813 188593 536049 188829
rect 535813 188273 536049 188509
rect 551952 188593 552188 188829
rect 551952 188273 552188 188509
rect 557882 188593 558118 188829
rect 557882 188273 558118 188509
rect 563813 188593 564049 188829
rect 563813 188273 564049 188509
rect 573526 188593 573762 188829
rect 573846 188593 574082 188829
rect 573526 188273 573762 188509
rect 573846 188273 574082 188509
rect 22916 185218 23152 185454
rect 22916 184898 23152 185134
rect 28847 185218 29083 185454
rect 28847 184898 29083 185134
rect 50916 185218 51152 185454
rect 50916 184898 51152 185134
rect 56847 185218 57083 185454
rect 56847 184898 57083 185134
rect 78916 185218 79152 185454
rect 78916 184898 79152 185134
rect 84847 185218 85083 185454
rect 84847 184898 85083 185134
rect 106916 185218 107152 185454
rect 106916 184898 107152 185134
rect 112847 185218 113083 185454
rect 112847 184898 113083 185134
rect 134916 185218 135152 185454
rect 134916 184898 135152 185134
rect 140847 185218 141083 185454
rect 140847 184898 141083 185134
rect 162916 185218 163152 185454
rect 162916 184898 163152 185134
rect 168847 185218 169083 185454
rect 168847 184898 169083 185134
rect 190916 185218 191152 185454
rect 190916 184898 191152 185134
rect 196847 185218 197083 185454
rect 196847 184898 197083 185134
rect 218916 185218 219152 185454
rect 218916 184898 219152 185134
rect 224847 185218 225083 185454
rect 224847 184898 225083 185134
rect 246916 185218 247152 185454
rect 246916 184898 247152 185134
rect 252847 185218 253083 185454
rect 252847 184898 253083 185134
rect 274916 185218 275152 185454
rect 274916 184898 275152 185134
rect 280847 185218 281083 185454
rect 280847 184898 281083 185134
rect 302916 185218 303152 185454
rect 302916 184898 303152 185134
rect 308847 185218 309083 185454
rect 308847 184898 309083 185134
rect 330916 185218 331152 185454
rect 330916 184898 331152 185134
rect 336847 185218 337083 185454
rect 336847 184898 337083 185134
rect 358916 185218 359152 185454
rect 358916 184898 359152 185134
rect 364847 185218 365083 185454
rect 364847 184898 365083 185134
rect 386916 185218 387152 185454
rect 386916 184898 387152 185134
rect 392847 185218 393083 185454
rect 392847 184898 393083 185134
rect 414916 185218 415152 185454
rect 414916 184898 415152 185134
rect 420847 185218 421083 185454
rect 420847 184898 421083 185134
rect 442916 185218 443152 185454
rect 442916 184898 443152 185134
rect 448847 185218 449083 185454
rect 448847 184898 449083 185134
rect 470916 185218 471152 185454
rect 470916 184898 471152 185134
rect 476847 185218 477083 185454
rect 476847 184898 477083 185134
rect 498916 185218 499152 185454
rect 498916 184898 499152 185134
rect 504847 185218 505083 185454
rect 504847 184898 505083 185134
rect 526916 185218 527152 185454
rect 526916 184898 527152 185134
rect 532847 185218 533083 185454
rect 532847 184898 533083 185134
rect 554916 185218 555152 185454
rect 554916 184898 555152 185134
rect 560847 185218 561083 185454
rect 560847 184898 561083 185134
rect -1974 161593 -1738 161829
rect -1654 161593 -1418 161829
rect -1974 161273 -1738 161509
rect -1654 161273 -1418 161509
rect 19952 161593 20188 161829
rect 19952 161273 20188 161509
rect 25882 161593 26118 161829
rect 25882 161273 26118 161509
rect 31813 161593 32049 161829
rect 31813 161273 32049 161509
rect 47952 161593 48188 161829
rect 47952 161273 48188 161509
rect 53882 161593 54118 161829
rect 53882 161273 54118 161509
rect 59813 161593 60049 161829
rect 59813 161273 60049 161509
rect 75952 161593 76188 161829
rect 75952 161273 76188 161509
rect 81882 161593 82118 161829
rect 81882 161273 82118 161509
rect 87813 161593 88049 161829
rect 87813 161273 88049 161509
rect 103952 161593 104188 161829
rect 103952 161273 104188 161509
rect 109882 161593 110118 161829
rect 109882 161273 110118 161509
rect 115813 161593 116049 161829
rect 115813 161273 116049 161509
rect 131952 161593 132188 161829
rect 131952 161273 132188 161509
rect 137882 161593 138118 161829
rect 137882 161273 138118 161509
rect 143813 161593 144049 161829
rect 143813 161273 144049 161509
rect 159952 161593 160188 161829
rect 159952 161273 160188 161509
rect 165882 161593 166118 161829
rect 165882 161273 166118 161509
rect 171813 161593 172049 161829
rect 171813 161273 172049 161509
rect 187952 161593 188188 161829
rect 187952 161273 188188 161509
rect 193882 161593 194118 161829
rect 193882 161273 194118 161509
rect 199813 161593 200049 161829
rect 199813 161273 200049 161509
rect 215952 161593 216188 161829
rect 215952 161273 216188 161509
rect 221882 161593 222118 161829
rect 221882 161273 222118 161509
rect 227813 161593 228049 161829
rect 227813 161273 228049 161509
rect 243952 161593 244188 161829
rect 243952 161273 244188 161509
rect 249882 161593 250118 161829
rect 249882 161273 250118 161509
rect 255813 161593 256049 161829
rect 255813 161273 256049 161509
rect 271952 161593 272188 161829
rect 271952 161273 272188 161509
rect 277882 161593 278118 161829
rect 277882 161273 278118 161509
rect 283813 161593 284049 161829
rect 283813 161273 284049 161509
rect 299952 161593 300188 161829
rect 299952 161273 300188 161509
rect 305882 161593 306118 161829
rect 305882 161273 306118 161509
rect 311813 161593 312049 161829
rect 311813 161273 312049 161509
rect 327952 161593 328188 161829
rect 327952 161273 328188 161509
rect 333882 161593 334118 161829
rect 333882 161273 334118 161509
rect 339813 161593 340049 161829
rect 339813 161273 340049 161509
rect 355952 161593 356188 161829
rect 355952 161273 356188 161509
rect 361882 161593 362118 161829
rect 361882 161273 362118 161509
rect 367813 161593 368049 161829
rect 367813 161273 368049 161509
rect 383952 161593 384188 161829
rect 383952 161273 384188 161509
rect 389882 161593 390118 161829
rect 389882 161273 390118 161509
rect 395813 161593 396049 161829
rect 395813 161273 396049 161509
rect 411952 161593 412188 161829
rect 411952 161273 412188 161509
rect 417882 161593 418118 161829
rect 417882 161273 418118 161509
rect 423813 161593 424049 161829
rect 423813 161273 424049 161509
rect 439952 161593 440188 161829
rect 439952 161273 440188 161509
rect 445882 161593 446118 161829
rect 445882 161273 446118 161509
rect 451813 161593 452049 161829
rect 451813 161273 452049 161509
rect 467952 161593 468188 161829
rect 467952 161273 468188 161509
rect 473882 161593 474118 161829
rect 473882 161273 474118 161509
rect 479813 161593 480049 161829
rect 479813 161273 480049 161509
rect 495952 161593 496188 161829
rect 495952 161273 496188 161509
rect 501882 161593 502118 161829
rect 501882 161273 502118 161509
rect 507813 161593 508049 161829
rect 507813 161273 508049 161509
rect 523952 161593 524188 161829
rect 523952 161273 524188 161509
rect 529882 161593 530118 161829
rect 529882 161273 530118 161509
rect 535813 161593 536049 161829
rect 535813 161273 536049 161509
rect 551952 161593 552188 161829
rect 551952 161273 552188 161509
rect 557882 161593 558118 161829
rect 557882 161273 558118 161509
rect 563813 161593 564049 161829
rect 563813 161273 564049 161509
rect 573526 161593 573762 161829
rect 573846 161593 574082 161829
rect 573526 161273 573762 161509
rect 573846 161273 574082 161509
rect 22916 158218 23152 158454
rect 22916 157898 23152 158134
rect 28847 158218 29083 158454
rect 28847 157898 29083 158134
rect 50916 158218 51152 158454
rect 50916 157898 51152 158134
rect 56847 158218 57083 158454
rect 56847 157898 57083 158134
rect 78916 158218 79152 158454
rect 78916 157898 79152 158134
rect 84847 158218 85083 158454
rect 84847 157898 85083 158134
rect 106916 158218 107152 158454
rect 106916 157898 107152 158134
rect 112847 158218 113083 158454
rect 112847 157898 113083 158134
rect 134916 158218 135152 158454
rect 134916 157898 135152 158134
rect 140847 158218 141083 158454
rect 140847 157898 141083 158134
rect 162916 158218 163152 158454
rect 162916 157898 163152 158134
rect 168847 158218 169083 158454
rect 168847 157898 169083 158134
rect 190916 158218 191152 158454
rect 190916 157898 191152 158134
rect 196847 158218 197083 158454
rect 196847 157898 197083 158134
rect 218916 158218 219152 158454
rect 218916 157898 219152 158134
rect 224847 158218 225083 158454
rect 224847 157898 225083 158134
rect 246916 158218 247152 158454
rect 246916 157898 247152 158134
rect 252847 158218 253083 158454
rect 252847 157898 253083 158134
rect 274916 158218 275152 158454
rect 274916 157898 275152 158134
rect 280847 158218 281083 158454
rect 280847 157898 281083 158134
rect 302916 158218 303152 158454
rect 302916 157898 303152 158134
rect 308847 158218 309083 158454
rect 308847 157898 309083 158134
rect 330916 158218 331152 158454
rect 330916 157898 331152 158134
rect 336847 158218 337083 158454
rect 336847 157898 337083 158134
rect 358916 158218 359152 158454
rect 358916 157898 359152 158134
rect 364847 158218 365083 158454
rect 364847 157898 365083 158134
rect 386916 158218 387152 158454
rect 386916 157898 387152 158134
rect 392847 158218 393083 158454
rect 392847 157898 393083 158134
rect 414916 158218 415152 158454
rect 414916 157898 415152 158134
rect 420847 158218 421083 158454
rect 420847 157898 421083 158134
rect 442916 158218 443152 158454
rect 442916 157898 443152 158134
rect 448847 158218 449083 158454
rect 448847 157898 449083 158134
rect 470916 158218 471152 158454
rect 470916 157898 471152 158134
rect 476847 158218 477083 158454
rect 476847 157898 477083 158134
rect 498916 158218 499152 158454
rect 498916 157898 499152 158134
rect 504847 158218 505083 158454
rect 504847 157898 505083 158134
rect 526916 158218 527152 158454
rect 526916 157898 527152 158134
rect 532847 158218 533083 158454
rect 532847 157898 533083 158134
rect 554916 158218 555152 158454
rect 554916 157898 555152 158134
rect 560847 158218 561083 158454
rect 560847 157898 561083 158134
rect -1974 134593 -1738 134829
rect -1654 134593 -1418 134829
rect -1974 134273 -1738 134509
rect -1654 134273 -1418 134509
rect 19952 134593 20188 134829
rect 19952 134273 20188 134509
rect 25882 134593 26118 134829
rect 25882 134273 26118 134509
rect 31813 134593 32049 134829
rect 31813 134273 32049 134509
rect 47952 134593 48188 134829
rect 47952 134273 48188 134509
rect 53882 134593 54118 134829
rect 53882 134273 54118 134509
rect 59813 134593 60049 134829
rect 59813 134273 60049 134509
rect 75952 134593 76188 134829
rect 75952 134273 76188 134509
rect 81882 134593 82118 134829
rect 81882 134273 82118 134509
rect 87813 134593 88049 134829
rect 87813 134273 88049 134509
rect 103952 134593 104188 134829
rect 103952 134273 104188 134509
rect 109882 134593 110118 134829
rect 109882 134273 110118 134509
rect 115813 134593 116049 134829
rect 115813 134273 116049 134509
rect 131952 134593 132188 134829
rect 131952 134273 132188 134509
rect 137882 134593 138118 134829
rect 137882 134273 138118 134509
rect 143813 134593 144049 134829
rect 143813 134273 144049 134509
rect 159952 134593 160188 134829
rect 159952 134273 160188 134509
rect 165882 134593 166118 134829
rect 165882 134273 166118 134509
rect 171813 134593 172049 134829
rect 171813 134273 172049 134509
rect 187952 134593 188188 134829
rect 187952 134273 188188 134509
rect 193882 134593 194118 134829
rect 193882 134273 194118 134509
rect 199813 134593 200049 134829
rect 199813 134273 200049 134509
rect 215952 134593 216188 134829
rect 215952 134273 216188 134509
rect 221882 134593 222118 134829
rect 221882 134273 222118 134509
rect 227813 134593 228049 134829
rect 227813 134273 228049 134509
rect 243952 134593 244188 134829
rect 243952 134273 244188 134509
rect 249882 134593 250118 134829
rect 249882 134273 250118 134509
rect 255813 134593 256049 134829
rect 255813 134273 256049 134509
rect 271952 134593 272188 134829
rect 271952 134273 272188 134509
rect 277882 134593 278118 134829
rect 277882 134273 278118 134509
rect 283813 134593 284049 134829
rect 283813 134273 284049 134509
rect 299952 134593 300188 134829
rect 299952 134273 300188 134509
rect 305882 134593 306118 134829
rect 305882 134273 306118 134509
rect 311813 134593 312049 134829
rect 311813 134273 312049 134509
rect 327952 134593 328188 134829
rect 327952 134273 328188 134509
rect 333882 134593 334118 134829
rect 333882 134273 334118 134509
rect 339813 134593 340049 134829
rect 339813 134273 340049 134509
rect 355952 134593 356188 134829
rect 355952 134273 356188 134509
rect 361882 134593 362118 134829
rect 361882 134273 362118 134509
rect 367813 134593 368049 134829
rect 367813 134273 368049 134509
rect 383952 134593 384188 134829
rect 383952 134273 384188 134509
rect 389882 134593 390118 134829
rect 389882 134273 390118 134509
rect 395813 134593 396049 134829
rect 395813 134273 396049 134509
rect 411952 134593 412188 134829
rect 411952 134273 412188 134509
rect 417882 134593 418118 134829
rect 417882 134273 418118 134509
rect 423813 134593 424049 134829
rect 423813 134273 424049 134509
rect 439952 134593 440188 134829
rect 439952 134273 440188 134509
rect 445882 134593 446118 134829
rect 445882 134273 446118 134509
rect 451813 134593 452049 134829
rect 451813 134273 452049 134509
rect 467952 134593 468188 134829
rect 467952 134273 468188 134509
rect 473882 134593 474118 134829
rect 473882 134273 474118 134509
rect 479813 134593 480049 134829
rect 479813 134273 480049 134509
rect 495952 134593 496188 134829
rect 495952 134273 496188 134509
rect 501882 134593 502118 134829
rect 501882 134273 502118 134509
rect 507813 134593 508049 134829
rect 507813 134273 508049 134509
rect 523952 134593 524188 134829
rect 523952 134273 524188 134509
rect 529882 134593 530118 134829
rect 529882 134273 530118 134509
rect 535813 134593 536049 134829
rect 535813 134273 536049 134509
rect 551952 134593 552188 134829
rect 551952 134273 552188 134509
rect 557882 134593 558118 134829
rect 557882 134273 558118 134509
rect 563813 134593 564049 134829
rect 563813 134273 564049 134509
rect 573526 134593 573762 134829
rect 573846 134593 574082 134829
rect 573526 134273 573762 134509
rect 573846 134273 574082 134509
rect 22916 131218 23152 131454
rect 22916 130898 23152 131134
rect 28847 131218 29083 131454
rect 28847 130898 29083 131134
rect 50916 131218 51152 131454
rect 50916 130898 51152 131134
rect 56847 131218 57083 131454
rect 56847 130898 57083 131134
rect 78916 131218 79152 131454
rect 78916 130898 79152 131134
rect 84847 131218 85083 131454
rect 84847 130898 85083 131134
rect 106916 131218 107152 131454
rect 106916 130898 107152 131134
rect 112847 131218 113083 131454
rect 112847 130898 113083 131134
rect 134916 131218 135152 131454
rect 134916 130898 135152 131134
rect 140847 131218 141083 131454
rect 140847 130898 141083 131134
rect 162916 131218 163152 131454
rect 162916 130898 163152 131134
rect 168847 131218 169083 131454
rect 168847 130898 169083 131134
rect 190916 131218 191152 131454
rect 190916 130898 191152 131134
rect 196847 131218 197083 131454
rect 196847 130898 197083 131134
rect 218916 131218 219152 131454
rect 218916 130898 219152 131134
rect 224847 131218 225083 131454
rect 224847 130898 225083 131134
rect 246916 131218 247152 131454
rect 246916 130898 247152 131134
rect 252847 131218 253083 131454
rect 252847 130898 253083 131134
rect 274916 131218 275152 131454
rect 274916 130898 275152 131134
rect 280847 131218 281083 131454
rect 280847 130898 281083 131134
rect 302916 131218 303152 131454
rect 302916 130898 303152 131134
rect 308847 131218 309083 131454
rect 308847 130898 309083 131134
rect 330916 131218 331152 131454
rect 330916 130898 331152 131134
rect 336847 131218 337083 131454
rect 336847 130898 337083 131134
rect 358916 131218 359152 131454
rect 358916 130898 359152 131134
rect 364847 131218 365083 131454
rect 364847 130898 365083 131134
rect 386916 131218 387152 131454
rect 386916 130898 387152 131134
rect 392847 131218 393083 131454
rect 392847 130898 393083 131134
rect 414916 131218 415152 131454
rect 414916 130898 415152 131134
rect 420847 131218 421083 131454
rect 420847 130898 421083 131134
rect 442916 131218 443152 131454
rect 442916 130898 443152 131134
rect 448847 131218 449083 131454
rect 448847 130898 449083 131134
rect 470916 131218 471152 131454
rect 470916 130898 471152 131134
rect 476847 131218 477083 131454
rect 476847 130898 477083 131134
rect 498916 131218 499152 131454
rect 498916 130898 499152 131134
rect 504847 131218 505083 131454
rect 504847 130898 505083 131134
rect 526916 131218 527152 131454
rect 526916 130898 527152 131134
rect 532847 131218 533083 131454
rect 532847 130898 533083 131134
rect 554916 131218 555152 131454
rect 554916 130898 555152 131134
rect 560847 131218 561083 131454
rect 560847 130898 561083 131134
rect -1974 107593 -1738 107829
rect -1654 107593 -1418 107829
rect -1974 107273 -1738 107509
rect -1654 107273 -1418 107509
rect 19952 107593 20188 107829
rect 19952 107273 20188 107509
rect 25882 107593 26118 107829
rect 25882 107273 26118 107509
rect 31813 107593 32049 107829
rect 31813 107273 32049 107509
rect 47952 107593 48188 107829
rect 47952 107273 48188 107509
rect 53882 107593 54118 107829
rect 53882 107273 54118 107509
rect 59813 107593 60049 107829
rect 59813 107273 60049 107509
rect 75952 107593 76188 107829
rect 75952 107273 76188 107509
rect 81882 107593 82118 107829
rect 81882 107273 82118 107509
rect 87813 107593 88049 107829
rect 87813 107273 88049 107509
rect 103952 107593 104188 107829
rect 103952 107273 104188 107509
rect 109882 107593 110118 107829
rect 109882 107273 110118 107509
rect 115813 107593 116049 107829
rect 115813 107273 116049 107509
rect 131952 107593 132188 107829
rect 131952 107273 132188 107509
rect 137882 107593 138118 107829
rect 137882 107273 138118 107509
rect 143813 107593 144049 107829
rect 143813 107273 144049 107509
rect 159952 107593 160188 107829
rect 159952 107273 160188 107509
rect 165882 107593 166118 107829
rect 165882 107273 166118 107509
rect 171813 107593 172049 107829
rect 171813 107273 172049 107509
rect 187952 107593 188188 107829
rect 187952 107273 188188 107509
rect 193882 107593 194118 107829
rect 193882 107273 194118 107509
rect 199813 107593 200049 107829
rect 199813 107273 200049 107509
rect 215952 107593 216188 107829
rect 215952 107273 216188 107509
rect 221882 107593 222118 107829
rect 221882 107273 222118 107509
rect 227813 107593 228049 107829
rect 227813 107273 228049 107509
rect 243952 107593 244188 107829
rect 243952 107273 244188 107509
rect 249882 107593 250118 107829
rect 249882 107273 250118 107509
rect 255813 107593 256049 107829
rect 255813 107273 256049 107509
rect 271952 107593 272188 107829
rect 271952 107273 272188 107509
rect 277882 107593 278118 107829
rect 277882 107273 278118 107509
rect 283813 107593 284049 107829
rect 283813 107273 284049 107509
rect 299952 107593 300188 107829
rect 299952 107273 300188 107509
rect 305882 107593 306118 107829
rect 305882 107273 306118 107509
rect 311813 107593 312049 107829
rect 311813 107273 312049 107509
rect 327952 107593 328188 107829
rect 327952 107273 328188 107509
rect 333882 107593 334118 107829
rect 333882 107273 334118 107509
rect 339813 107593 340049 107829
rect 339813 107273 340049 107509
rect 355952 107593 356188 107829
rect 355952 107273 356188 107509
rect 361882 107593 362118 107829
rect 361882 107273 362118 107509
rect 367813 107593 368049 107829
rect 367813 107273 368049 107509
rect 383952 107593 384188 107829
rect 383952 107273 384188 107509
rect 389882 107593 390118 107829
rect 389882 107273 390118 107509
rect 395813 107593 396049 107829
rect 395813 107273 396049 107509
rect 411952 107593 412188 107829
rect 411952 107273 412188 107509
rect 417882 107593 418118 107829
rect 417882 107273 418118 107509
rect 423813 107593 424049 107829
rect 423813 107273 424049 107509
rect 439952 107593 440188 107829
rect 439952 107273 440188 107509
rect 445882 107593 446118 107829
rect 445882 107273 446118 107509
rect 451813 107593 452049 107829
rect 451813 107273 452049 107509
rect 467952 107593 468188 107829
rect 467952 107273 468188 107509
rect 473882 107593 474118 107829
rect 473882 107273 474118 107509
rect 479813 107593 480049 107829
rect 479813 107273 480049 107509
rect 495952 107593 496188 107829
rect 495952 107273 496188 107509
rect 501882 107593 502118 107829
rect 501882 107273 502118 107509
rect 507813 107593 508049 107829
rect 507813 107273 508049 107509
rect 523952 107593 524188 107829
rect 523952 107273 524188 107509
rect 529882 107593 530118 107829
rect 529882 107273 530118 107509
rect 535813 107593 536049 107829
rect 535813 107273 536049 107509
rect 551952 107593 552188 107829
rect 551952 107273 552188 107509
rect 557882 107593 558118 107829
rect 557882 107273 558118 107509
rect 563813 107593 564049 107829
rect 563813 107273 564049 107509
rect 573526 107593 573762 107829
rect 573846 107593 574082 107829
rect 573526 107273 573762 107509
rect 573846 107273 574082 107509
rect 22916 104218 23152 104454
rect 22916 103898 23152 104134
rect 28847 104218 29083 104454
rect 28847 103898 29083 104134
rect 50916 104218 51152 104454
rect 50916 103898 51152 104134
rect 56847 104218 57083 104454
rect 56847 103898 57083 104134
rect 78916 104218 79152 104454
rect 78916 103898 79152 104134
rect 84847 104218 85083 104454
rect 84847 103898 85083 104134
rect 106916 104218 107152 104454
rect 106916 103898 107152 104134
rect 112847 104218 113083 104454
rect 112847 103898 113083 104134
rect 134916 104218 135152 104454
rect 134916 103898 135152 104134
rect 140847 104218 141083 104454
rect 140847 103898 141083 104134
rect 162916 104218 163152 104454
rect 162916 103898 163152 104134
rect 168847 104218 169083 104454
rect 168847 103898 169083 104134
rect 190916 104218 191152 104454
rect 190916 103898 191152 104134
rect 196847 104218 197083 104454
rect 196847 103898 197083 104134
rect 218916 104218 219152 104454
rect 218916 103898 219152 104134
rect 224847 104218 225083 104454
rect 224847 103898 225083 104134
rect 246916 104218 247152 104454
rect 246916 103898 247152 104134
rect 252847 104218 253083 104454
rect 252847 103898 253083 104134
rect 274916 104218 275152 104454
rect 274916 103898 275152 104134
rect 280847 104218 281083 104454
rect 280847 103898 281083 104134
rect 302916 104218 303152 104454
rect 302916 103898 303152 104134
rect 308847 104218 309083 104454
rect 308847 103898 309083 104134
rect 330916 104218 331152 104454
rect 330916 103898 331152 104134
rect 336847 104218 337083 104454
rect 336847 103898 337083 104134
rect 358916 104218 359152 104454
rect 358916 103898 359152 104134
rect 364847 104218 365083 104454
rect 364847 103898 365083 104134
rect 386916 104218 387152 104454
rect 386916 103898 387152 104134
rect 392847 104218 393083 104454
rect 392847 103898 393083 104134
rect 414916 104218 415152 104454
rect 414916 103898 415152 104134
rect 420847 104218 421083 104454
rect 420847 103898 421083 104134
rect 442916 104218 443152 104454
rect 442916 103898 443152 104134
rect 448847 104218 449083 104454
rect 448847 103898 449083 104134
rect 470916 104218 471152 104454
rect 470916 103898 471152 104134
rect 476847 104218 477083 104454
rect 476847 103898 477083 104134
rect 498916 104218 499152 104454
rect 498916 103898 499152 104134
rect 504847 104218 505083 104454
rect 504847 103898 505083 104134
rect 526916 104218 527152 104454
rect 526916 103898 527152 104134
rect 532847 104218 533083 104454
rect 532847 103898 533083 104134
rect 554916 104218 555152 104454
rect 554916 103898 555152 104134
rect 560847 104218 561083 104454
rect 560847 103898 561083 104134
rect -1974 80593 -1738 80829
rect -1654 80593 -1418 80829
rect -1974 80273 -1738 80509
rect -1654 80273 -1418 80509
rect 19952 80593 20188 80829
rect 19952 80273 20188 80509
rect 25882 80593 26118 80829
rect 25882 80273 26118 80509
rect 31813 80593 32049 80829
rect 31813 80273 32049 80509
rect 47952 80593 48188 80829
rect 47952 80273 48188 80509
rect 53882 80593 54118 80829
rect 53882 80273 54118 80509
rect 59813 80593 60049 80829
rect 59813 80273 60049 80509
rect 75952 80593 76188 80829
rect 75952 80273 76188 80509
rect 81882 80593 82118 80829
rect 81882 80273 82118 80509
rect 87813 80593 88049 80829
rect 87813 80273 88049 80509
rect 103952 80593 104188 80829
rect 103952 80273 104188 80509
rect 109882 80593 110118 80829
rect 109882 80273 110118 80509
rect 115813 80593 116049 80829
rect 115813 80273 116049 80509
rect 131952 80593 132188 80829
rect 131952 80273 132188 80509
rect 137882 80593 138118 80829
rect 137882 80273 138118 80509
rect 143813 80593 144049 80829
rect 143813 80273 144049 80509
rect 159952 80593 160188 80829
rect 159952 80273 160188 80509
rect 165882 80593 166118 80829
rect 165882 80273 166118 80509
rect 171813 80593 172049 80829
rect 171813 80273 172049 80509
rect 187952 80593 188188 80829
rect 187952 80273 188188 80509
rect 193882 80593 194118 80829
rect 193882 80273 194118 80509
rect 199813 80593 200049 80829
rect 199813 80273 200049 80509
rect 215952 80593 216188 80829
rect 215952 80273 216188 80509
rect 221882 80593 222118 80829
rect 221882 80273 222118 80509
rect 227813 80593 228049 80829
rect 227813 80273 228049 80509
rect 243952 80593 244188 80829
rect 243952 80273 244188 80509
rect 249882 80593 250118 80829
rect 249882 80273 250118 80509
rect 255813 80593 256049 80829
rect 255813 80273 256049 80509
rect 271952 80593 272188 80829
rect 271952 80273 272188 80509
rect 277882 80593 278118 80829
rect 277882 80273 278118 80509
rect 283813 80593 284049 80829
rect 283813 80273 284049 80509
rect 299952 80593 300188 80829
rect 299952 80273 300188 80509
rect 305882 80593 306118 80829
rect 305882 80273 306118 80509
rect 311813 80593 312049 80829
rect 311813 80273 312049 80509
rect 327952 80593 328188 80829
rect 327952 80273 328188 80509
rect 333882 80593 334118 80829
rect 333882 80273 334118 80509
rect 339813 80593 340049 80829
rect 339813 80273 340049 80509
rect 355952 80593 356188 80829
rect 355952 80273 356188 80509
rect 361882 80593 362118 80829
rect 361882 80273 362118 80509
rect 367813 80593 368049 80829
rect 367813 80273 368049 80509
rect 383952 80593 384188 80829
rect 383952 80273 384188 80509
rect 389882 80593 390118 80829
rect 389882 80273 390118 80509
rect 395813 80593 396049 80829
rect 395813 80273 396049 80509
rect 411952 80593 412188 80829
rect 411952 80273 412188 80509
rect 417882 80593 418118 80829
rect 417882 80273 418118 80509
rect 423813 80593 424049 80829
rect 423813 80273 424049 80509
rect 439952 80593 440188 80829
rect 439952 80273 440188 80509
rect 445882 80593 446118 80829
rect 445882 80273 446118 80509
rect 451813 80593 452049 80829
rect 451813 80273 452049 80509
rect 467952 80593 468188 80829
rect 467952 80273 468188 80509
rect 473882 80593 474118 80829
rect 473882 80273 474118 80509
rect 479813 80593 480049 80829
rect 479813 80273 480049 80509
rect 495952 80593 496188 80829
rect 495952 80273 496188 80509
rect 501882 80593 502118 80829
rect 501882 80273 502118 80509
rect 507813 80593 508049 80829
rect 507813 80273 508049 80509
rect 523952 80593 524188 80829
rect 523952 80273 524188 80509
rect 529882 80593 530118 80829
rect 529882 80273 530118 80509
rect 535813 80593 536049 80829
rect 535813 80273 536049 80509
rect 551952 80593 552188 80829
rect 551952 80273 552188 80509
rect 557882 80593 558118 80829
rect 557882 80273 558118 80509
rect 563813 80593 564049 80829
rect 563813 80273 564049 80509
rect 573526 80593 573762 80829
rect 573846 80593 574082 80829
rect 573526 80273 573762 80509
rect 573846 80273 574082 80509
rect 22916 77218 23152 77454
rect 22916 76898 23152 77134
rect 28847 77218 29083 77454
rect 28847 76898 29083 77134
rect 50916 77218 51152 77454
rect 50916 76898 51152 77134
rect 56847 77218 57083 77454
rect 56847 76898 57083 77134
rect 78916 77218 79152 77454
rect 78916 76898 79152 77134
rect 84847 77218 85083 77454
rect 84847 76898 85083 77134
rect 106916 77218 107152 77454
rect 106916 76898 107152 77134
rect 112847 77218 113083 77454
rect 112847 76898 113083 77134
rect 134916 77218 135152 77454
rect 134916 76898 135152 77134
rect 140847 77218 141083 77454
rect 140847 76898 141083 77134
rect 162916 77218 163152 77454
rect 162916 76898 163152 77134
rect 168847 77218 169083 77454
rect 168847 76898 169083 77134
rect 190916 77218 191152 77454
rect 190916 76898 191152 77134
rect 196847 77218 197083 77454
rect 196847 76898 197083 77134
rect 218916 77218 219152 77454
rect 218916 76898 219152 77134
rect 224847 77218 225083 77454
rect 224847 76898 225083 77134
rect 246916 77218 247152 77454
rect 246916 76898 247152 77134
rect 252847 77218 253083 77454
rect 252847 76898 253083 77134
rect 274916 77218 275152 77454
rect 274916 76898 275152 77134
rect 280847 77218 281083 77454
rect 280847 76898 281083 77134
rect 302916 77218 303152 77454
rect 302916 76898 303152 77134
rect 308847 77218 309083 77454
rect 308847 76898 309083 77134
rect 330916 77218 331152 77454
rect 330916 76898 331152 77134
rect 336847 77218 337083 77454
rect 336847 76898 337083 77134
rect 358916 77218 359152 77454
rect 358916 76898 359152 77134
rect 364847 77218 365083 77454
rect 364847 76898 365083 77134
rect 386916 77218 387152 77454
rect 386916 76898 387152 77134
rect 392847 77218 393083 77454
rect 392847 76898 393083 77134
rect 414916 77218 415152 77454
rect 414916 76898 415152 77134
rect 420847 77218 421083 77454
rect 420847 76898 421083 77134
rect 442916 77218 443152 77454
rect 442916 76898 443152 77134
rect 448847 77218 449083 77454
rect 448847 76898 449083 77134
rect 470916 77218 471152 77454
rect 470916 76898 471152 77134
rect 476847 77218 477083 77454
rect 476847 76898 477083 77134
rect 498916 77218 499152 77454
rect 498916 76898 499152 77134
rect 504847 77218 505083 77454
rect 504847 76898 505083 77134
rect 526916 77218 527152 77454
rect 526916 76898 527152 77134
rect 532847 77218 533083 77454
rect 532847 76898 533083 77134
rect 554916 77218 555152 77454
rect 554916 76898 555152 77134
rect 560847 77218 561083 77454
rect 560847 76898 561083 77134
rect -1974 53593 -1738 53829
rect -1654 53593 -1418 53829
rect -1974 53273 -1738 53509
rect -1654 53273 -1418 53509
rect 19952 53593 20188 53829
rect 19952 53273 20188 53509
rect 25882 53593 26118 53829
rect 25882 53273 26118 53509
rect 31813 53593 32049 53829
rect 31813 53273 32049 53509
rect 47952 53593 48188 53829
rect 47952 53273 48188 53509
rect 53882 53593 54118 53829
rect 53882 53273 54118 53509
rect 59813 53593 60049 53829
rect 59813 53273 60049 53509
rect 75952 53593 76188 53829
rect 75952 53273 76188 53509
rect 81882 53593 82118 53829
rect 81882 53273 82118 53509
rect 87813 53593 88049 53829
rect 87813 53273 88049 53509
rect 103952 53593 104188 53829
rect 103952 53273 104188 53509
rect 109882 53593 110118 53829
rect 109882 53273 110118 53509
rect 115813 53593 116049 53829
rect 115813 53273 116049 53509
rect 131952 53593 132188 53829
rect 131952 53273 132188 53509
rect 137882 53593 138118 53829
rect 137882 53273 138118 53509
rect 143813 53593 144049 53829
rect 143813 53273 144049 53509
rect 159952 53593 160188 53829
rect 159952 53273 160188 53509
rect 165882 53593 166118 53829
rect 165882 53273 166118 53509
rect 171813 53593 172049 53829
rect 171813 53273 172049 53509
rect 187952 53593 188188 53829
rect 187952 53273 188188 53509
rect 193882 53593 194118 53829
rect 193882 53273 194118 53509
rect 199813 53593 200049 53829
rect 199813 53273 200049 53509
rect 215952 53593 216188 53829
rect 215952 53273 216188 53509
rect 221882 53593 222118 53829
rect 221882 53273 222118 53509
rect 227813 53593 228049 53829
rect 227813 53273 228049 53509
rect 243952 53593 244188 53829
rect 243952 53273 244188 53509
rect 249882 53593 250118 53829
rect 249882 53273 250118 53509
rect 255813 53593 256049 53829
rect 255813 53273 256049 53509
rect 271952 53593 272188 53829
rect 271952 53273 272188 53509
rect 277882 53593 278118 53829
rect 277882 53273 278118 53509
rect 283813 53593 284049 53829
rect 283813 53273 284049 53509
rect 299952 53593 300188 53829
rect 299952 53273 300188 53509
rect 305882 53593 306118 53829
rect 305882 53273 306118 53509
rect 311813 53593 312049 53829
rect 311813 53273 312049 53509
rect 327952 53593 328188 53829
rect 327952 53273 328188 53509
rect 333882 53593 334118 53829
rect 333882 53273 334118 53509
rect 339813 53593 340049 53829
rect 339813 53273 340049 53509
rect 355952 53593 356188 53829
rect 355952 53273 356188 53509
rect 361882 53593 362118 53829
rect 361882 53273 362118 53509
rect 367813 53593 368049 53829
rect 367813 53273 368049 53509
rect 383952 53593 384188 53829
rect 383952 53273 384188 53509
rect 389882 53593 390118 53829
rect 389882 53273 390118 53509
rect 395813 53593 396049 53829
rect 395813 53273 396049 53509
rect 411952 53593 412188 53829
rect 411952 53273 412188 53509
rect 417882 53593 418118 53829
rect 417882 53273 418118 53509
rect 423813 53593 424049 53829
rect 423813 53273 424049 53509
rect 439952 53593 440188 53829
rect 439952 53273 440188 53509
rect 445882 53593 446118 53829
rect 445882 53273 446118 53509
rect 451813 53593 452049 53829
rect 451813 53273 452049 53509
rect 467952 53593 468188 53829
rect 467952 53273 468188 53509
rect 473882 53593 474118 53829
rect 473882 53273 474118 53509
rect 479813 53593 480049 53829
rect 479813 53273 480049 53509
rect 495952 53593 496188 53829
rect 495952 53273 496188 53509
rect 501882 53593 502118 53829
rect 501882 53273 502118 53509
rect 507813 53593 508049 53829
rect 507813 53273 508049 53509
rect 523952 53593 524188 53829
rect 523952 53273 524188 53509
rect 529882 53593 530118 53829
rect 529882 53273 530118 53509
rect 535813 53593 536049 53829
rect 535813 53273 536049 53509
rect 551952 53593 552188 53829
rect 551952 53273 552188 53509
rect 557882 53593 558118 53829
rect 557882 53273 558118 53509
rect 563813 53593 564049 53829
rect 563813 53273 564049 53509
rect 573526 53593 573762 53829
rect 573846 53593 574082 53829
rect 573526 53273 573762 53509
rect 573846 53273 574082 53509
rect 22916 50218 23152 50454
rect 22916 49898 23152 50134
rect 28847 50218 29083 50454
rect 28847 49898 29083 50134
rect 50916 50218 51152 50454
rect 50916 49898 51152 50134
rect 56847 50218 57083 50454
rect 56847 49898 57083 50134
rect 78916 50218 79152 50454
rect 78916 49898 79152 50134
rect 84847 50218 85083 50454
rect 84847 49898 85083 50134
rect 106916 50218 107152 50454
rect 106916 49898 107152 50134
rect 112847 50218 113083 50454
rect 112847 49898 113083 50134
rect 134916 50218 135152 50454
rect 134916 49898 135152 50134
rect 140847 50218 141083 50454
rect 140847 49898 141083 50134
rect 162916 50218 163152 50454
rect 162916 49898 163152 50134
rect 168847 50218 169083 50454
rect 168847 49898 169083 50134
rect 190916 50218 191152 50454
rect 190916 49898 191152 50134
rect 196847 50218 197083 50454
rect 196847 49898 197083 50134
rect 218916 50218 219152 50454
rect 218916 49898 219152 50134
rect 224847 50218 225083 50454
rect 224847 49898 225083 50134
rect 246916 50218 247152 50454
rect 246916 49898 247152 50134
rect 252847 50218 253083 50454
rect 252847 49898 253083 50134
rect 274916 50218 275152 50454
rect 274916 49898 275152 50134
rect 280847 50218 281083 50454
rect 280847 49898 281083 50134
rect 302916 50218 303152 50454
rect 302916 49898 303152 50134
rect 308847 50218 309083 50454
rect 308847 49898 309083 50134
rect 330916 50218 331152 50454
rect 330916 49898 331152 50134
rect 336847 50218 337083 50454
rect 336847 49898 337083 50134
rect 358916 50218 359152 50454
rect 358916 49898 359152 50134
rect 364847 50218 365083 50454
rect 364847 49898 365083 50134
rect 386916 50218 387152 50454
rect 386916 49898 387152 50134
rect 392847 50218 393083 50454
rect 392847 49898 393083 50134
rect 414916 50218 415152 50454
rect 414916 49898 415152 50134
rect 420847 50218 421083 50454
rect 420847 49898 421083 50134
rect 442916 50218 443152 50454
rect 442916 49898 443152 50134
rect 448847 50218 449083 50454
rect 448847 49898 449083 50134
rect 470916 50218 471152 50454
rect 470916 49898 471152 50134
rect 476847 50218 477083 50454
rect 476847 49898 477083 50134
rect 498916 50218 499152 50454
rect 498916 49898 499152 50134
rect 504847 50218 505083 50454
rect 504847 49898 505083 50134
rect 526916 50218 527152 50454
rect 526916 49898 527152 50134
rect 532847 50218 533083 50454
rect 532847 49898 533083 50134
rect 554916 50218 555152 50454
rect 554916 49898 555152 50134
rect 560847 50218 561083 50454
rect 560847 49898 561083 50134
rect -1974 26593 -1738 26829
rect -1654 26593 -1418 26829
rect -1974 26273 -1738 26509
rect -1654 26273 -1418 26509
rect 24284 26593 24520 26829
rect 24284 26273 24520 26509
rect 38882 26593 39118 26829
rect 38882 26273 39118 26509
rect 53479 26593 53715 26829
rect 53479 26273 53715 26509
rect 31584 23218 31820 23454
rect 31584 22898 31820 23134
rect 46181 23218 46417 23454
rect 46181 22898 46417 23134
rect 75952 26593 76188 26829
rect 75952 26273 76188 26509
rect 81882 26593 82118 26829
rect 81882 26273 82118 26509
rect 87813 26593 88049 26829
rect 87813 26273 88049 26509
rect 103952 26593 104188 26829
rect 103952 26273 104188 26509
rect 109882 26593 110118 26829
rect 109882 26273 110118 26509
rect 115813 26593 116049 26829
rect 115813 26273 116049 26509
rect 131952 26593 132188 26829
rect 131952 26273 132188 26509
rect 137882 26593 138118 26829
rect 137882 26273 138118 26509
rect 143813 26593 144049 26829
rect 143813 26273 144049 26509
rect 159952 26593 160188 26829
rect 159952 26273 160188 26509
rect 165882 26593 166118 26829
rect 165882 26273 166118 26509
rect 171813 26593 172049 26829
rect 171813 26273 172049 26509
rect 187952 26593 188188 26829
rect 187952 26273 188188 26509
rect 193882 26593 194118 26829
rect 193882 26273 194118 26509
rect 199813 26593 200049 26829
rect 199813 26273 200049 26509
rect 215952 26593 216188 26829
rect 215952 26273 216188 26509
rect 221882 26593 222118 26829
rect 221882 26273 222118 26509
rect 227813 26593 228049 26829
rect 227813 26273 228049 26509
rect 243952 26593 244188 26829
rect 243952 26273 244188 26509
rect 249882 26593 250118 26829
rect 249882 26273 250118 26509
rect 255813 26593 256049 26829
rect 255813 26273 256049 26509
rect 271952 26593 272188 26829
rect 271952 26273 272188 26509
rect 277882 26593 278118 26829
rect 277882 26273 278118 26509
rect 283813 26593 284049 26829
rect 283813 26273 284049 26509
rect 299952 26593 300188 26829
rect 299952 26273 300188 26509
rect 305882 26593 306118 26829
rect 305882 26273 306118 26509
rect 311813 26593 312049 26829
rect 311813 26273 312049 26509
rect 327952 26593 328188 26829
rect 327952 26273 328188 26509
rect 333882 26593 334118 26829
rect 333882 26273 334118 26509
rect 339813 26593 340049 26829
rect 339813 26273 340049 26509
rect 355952 26593 356188 26829
rect 355952 26273 356188 26509
rect 361882 26593 362118 26829
rect 361882 26273 362118 26509
rect 367813 26593 368049 26829
rect 367813 26273 368049 26509
rect 383952 26593 384188 26829
rect 383952 26273 384188 26509
rect 389882 26593 390118 26829
rect 389882 26273 390118 26509
rect 395813 26593 396049 26829
rect 395813 26273 396049 26509
rect 411952 26593 412188 26829
rect 411952 26273 412188 26509
rect 417882 26593 418118 26829
rect 417882 26273 418118 26509
rect 423813 26593 424049 26829
rect 423813 26273 424049 26509
rect 439952 26593 440188 26829
rect 439952 26273 440188 26509
rect 445882 26593 446118 26829
rect 445882 26273 446118 26509
rect 451813 26593 452049 26829
rect 451813 26273 452049 26509
rect 467952 26593 468188 26829
rect 467952 26273 468188 26509
rect 473882 26593 474118 26829
rect 473882 26273 474118 26509
rect 479813 26593 480049 26829
rect 479813 26273 480049 26509
rect 495952 26593 496188 26829
rect 495952 26273 496188 26509
rect 501882 26593 502118 26829
rect 501882 26273 502118 26509
rect 507813 26593 508049 26829
rect 507813 26273 508049 26509
rect 523952 26593 524188 26829
rect 523952 26273 524188 26509
rect 529882 26593 530118 26829
rect 529882 26273 530118 26509
rect 535813 26593 536049 26829
rect 535813 26273 536049 26509
rect 551952 26593 552188 26829
rect 551952 26273 552188 26509
rect 557882 26593 558118 26829
rect 557882 26273 558118 26509
rect 563813 26593 564049 26829
rect 563813 26273 564049 26509
rect 573526 26593 573762 26829
rect 573846 26593 574082 26829
rect 573526 26273 573762 26509
rect 573846 26273 574082 26509
rect 66026 23218 66262 23454
rect 66346 23218 66582 23454
rect 66026 22898 66262 23134
rect 66346 22898 66582 23134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 78916 23218 79152 23454
rect 78916 22898 79152 23134
rect 84847 23218 85083 23454
rect 84847 22898 85083 23134
rect 106916 23218 107152 23454
rect 106916 22898 107152 23134
rect 112847 23218 113083 23454
rect 112847 22898 113083 23134
rect 134916 23218 135152 23454
rect 134916 22898 135152 23134
rect 140847 23218 141083 23454
rect 140847 22898 141083 23134
rect 162916 23218 163152 23454
rect 162916 22898 163152 23134
rect 168847 23218 169083 23454
rect 168847 22898 169083 23134
rect 190916 23218 191152 23454
rect 190916 22898 191152 23134
rect 196847 23218 197083 23454
rect 196847 22898 197083 23134
rect 218916 23218 219152 23454
rect 218916 22898 219152 23134
rect 224847 23218 225083 23454
rect 224847 22898 225083 23134
rect 246916 23218 247152 23454
rect 246916 22898 247152 23134
rect 252847 23218 253083 23454
rect 252847 22898 253083 23134
rect 274916 23218 275152 23454
rect 274916 22898 275152 23134
rect 280847 23218 281083 23454
rect 280847 22898 281083 23134
rect 302916 23218 303152 23454
rect 302916 22898 303152 23134
rect 308847 23218 309083 23454
rect 308847 22898 309083 23134
rect 330916 23218 331152 23454
rect 330916 22898 331152 23134
rect 336847 23218 337083 23454
rect 336847 22898 337083 23134
rect 358916 23218 359152 23454
rect 358916 22898 359152 23134
rect 364847 23218 365083 23454
rect 364847 22898 365083 23134
rect 386916 23218 387152 23454
rect 386916 22898 387152 23134
rect 392847 23218 393083 23454
rect 392847 22898 393083 23134
rect 414916 23218 415152 23454
rect 414916 22898 415152 23134
rect 420847 23218 421083 23454
rect 420847 22898 421083 23134
rect 442916 23218 443152 23454
rect 442916 22898 443152 23134
rect 448847 23218 449083 23454
rect 448847 22898 449083 23134
rect 470916 23218 471152 23454
rect 470916 22898 471152 23134
rect 476847 23218 477083 23454
rect 476847 22898 477083 23134
rect 498916 23218 499152 23454
rect 498916 22898 499152 23134
rect 504847 23218 505083 23454
rect 504847 22898 505083 23134
rect 526916 23218 527152 23454
rect 526916 22898 527152 23134
rect 532847 23218 533083 23454
rect 532847 22898 533083 23134
rect 554916 23218 555152 23454
rect 554916 22898 555152 23134
rect 560847 23218 561083 23454
rect 560847 22898 561083 23134
rect 66026 -1542 66262 -1306
rect 66346 -1542 66582 -1306
rect 66026 -1862 66262 -1626
rect 66346 -1862 66582 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 573526 -582 573762 -346
rect 573846 -582 574082 -346
rect 573526 -902 573762 -666
rect 573846 -902 574082 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 701593 585578 701829
rect 585662 701593 585898 701829
rect 585342 701273 585578 701509
rect 585662 701273 585898 701509
rect 585342 674593 585578 674829
rect 585662 674593 585898 674829
rect 585342 674273 585578 674509
rect 585662 674273 585898 674509
rect 585342 647593 585578 647829
rect 585662 647593 585898 647829
rect 585342 647273 585578 647509
rect 585662 647273 585898 647509
rect 585342 620593 585578 620829
rect 585662 620593 585898 620829
rect 585342 620273 585578 620509
rect 585662 620273 585898 620509
rect 585342 593593 585578 593829
rect 585662 593593 585898 593829
rect 585342 593273 585578 593509
rect 585662 593273 585898 593509
rect 585342 566593 585578 566829
rect 585662 566593 585898 566829
rect 585342 566273 585578 566509
rect 585662 566273 585898 566509
rect 585342 539593 585578 539829
rect 585662 539593 585898 539829
rect 585342 539273 585578 539509
rect 585662 539273 585898 539509
rect 585342 512593 585578 512829
rect 585662 512593 585898 512829
rect 585342 512273 585578 512509
rect 585662 512273 585898 512509
rect 585342 485593 585578 485829
rect 585662 485593 585898 485829
rect 585342 485273 585578 485509
rect 585662 485273 585898 485509
rect 585342 458593 585578 458829
rect 585662 458593 585898 458829
rect 585342 458273 585578 458509
rect 585662 458273 585898 458509
rect 585342 431593 585578 431829
rect 585662 431593 585898 431829
rect 585342 431273 585578 431509
rect 585662 431273 585898 431509
rect 585342 404593 585578 404829
rect 585662 404593 585898 404829
rect 585342 404273 585578 404509
rect 585662 404273 585898 404509
rect 585342 377593 585578 377829
rect 585662 377593 585898 377829
rect 585342 377273 585578 377509
rect 585662 377273 585898 377509
rect 585342 350593 585578 350829
rect 585662 350593 585898 350829
rect 585342 350273 585578 350509
rect 585662 350273 585898 350509
rect 585342 323593 585578 323829
rect 585662 323593 585898 323829
rect 585342 323273 585578 323509
rect 585662 323273 585898 323509
rect 585342 296593 585578 296829
rect 585662 296593 585898 296829
rect 585342 296273 585578 296509
rect 585662 296273 585898 296509
rect 585342 269593 585578 269829
rect 585662 269593 585898 269829
rect 585342 269273 585578 269509
rect 585662 269273 585898 269509
rect 585342 242593 585578 242829
rect 585662 242593 585898 242829
rect 585342 242273 585578 242509
rect 585662 242273 585898 242509
rect 585342 215593 585578 215829
rect 585662 215593 585898 215829
rect 585342 215273 585578 215509
rect 585662 215273 585898 215509
rect 585342 188593 585578 188829
rect 585662 188593 585898 188829
rect 585342 188273 585578 188509
rect 585662 188273 585898 188509
rect 585342 161593 585578 161829
rect 585662 161593 585898 161829
rect 585342 161273 585578 161509
rect 585662 161273 585898 161509
rect 585342 134593 585578 134829
rect 585662 134593 585898 134829
rect 585342 134273 585578 134509
rect 585662 134273 585898 134509
rect 585342 107593 585578 107829
rect 585662 107593 585898 107829
rect 585342 107273 585578 107509
rect 585662 107273 585898 107509
rect 585342 80593 585578 80829
rect 585662 80593 585898 80829
rect 585342 80273 585578 80509
rect 585662 80273 585898 80509
rect 585342 53593 585578 53829
rect 585662 53593 585898 53829
rect 585342 53273 585578 53509
rect 585662 53273 585898 53509
rect 585342 26593 585578 26829
rect 585662 26593 585898 26829
rect 585342 26273 585578 26509
rect 585662 26273 585898 26509
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 698218 586538 698454
rect 586622 698218 586858 698454
rect 586302 697898 586538 698134
rect 586622 697898 586858 698134
rect 586302 671218 586538 671454
rect 586622 671218 586858 671454
rect 586302 670898 586538 671134
rect 586622 670898 586858 671134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 617218 586538 617454
rect 586622 617218 586858 617454
rect 586302 616898 586538 617134
rect 586622 616898 586858 617134
rect 586302 590218 586538 590454
rect 586622 590218 586858 590454
rect 586302 589898 586538 590134
rect 586622 589898 586858 590134
rect 586302 563218 586538 563454
rect 586622 563218 586858 563454
rect 586302 562898 586538 563134
rect 586622 562898 586858 563134
rect 586302 536218 586538 536454
rect 586622 536218 586858 536454
rect 586302 535898 586538 536134
rect 586622 535898 586858 536134
rect 586302 509218 586538 509454
rect 586622 509218 586858 509454
rect 586302 508898 586538 509134
rect 586622 508898 586858 509134
rect 586302 482218 586538 482454
rect 586622 482218 586858 482454
rect 586302 481898 586538 482134
rect 586622 481898 586858 482134
rect 586302 455218 586538 455454
rect 586622 455218 586858 455454
rect 586302 454898 586538 455134
rect 586622 454898 586858 455134
rect 586302 428218 586538 428454
rect 586622 428218 586858 428454
rect 586302 427898 586538 428134
rect 586622 427898 586858 428134
rect 586302 401218 586538 401454
rect 586622 401218 586858 401454
rect 586302 400898 586538 401134
rect 586622 400898 586858 401134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 347218 586538 347454
rect 586622 347218 586858 347454
rect 586302 346898 586538 347134
rect 586622 346898 586858 347134
rect 586302 320218 586538 320454
rect 586622 320218 586858 320454
rect 586302 319898 586538 320134
rect 586622 319898 586858 320134
rect 586302 293218 586538 293454
rect 586622 293218 586858 293454
rect 586302 292898 586538 293134
rect 586622 292898 586858 293134
rect 586302 266218 586538 266454
rect 586622 266218 586858 266454
rect 586302 265898 586538 266134
rect 586622 265898 586858 266134
rect 586302 239218 586538 239454
rect 586622 239218 586858 239454
rect 586302 238898 586538 239134
rect 586622 238898 586858 239134
rect 586302 212218 586538 212454
rect 586622 212218 586858 212454
rect 586302 211898 586538 212134
rect 586622 211898 586858 212134
rect 586302 185218 586538 185454
rect 586622 185218 586858 185454
rect 586302 184898 586538 185134
rect 586622 184898 586858 185134
rect 586302 158218 586538 158454
rect 586622 158218 586858 158454
rect 586302 157898 586538 158134
rect 586622 157898 586858 158134
rect 586302 131218 586538 131454
rect 586622 131218 586858 131454
rect 586302 130898 586538 131134
rect 586622 130898 586858 131134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 77218 586538 77454
rect 586622 77218 586858 77454
rect 586302 76898 586538 77134
rect 586622 76898 586858 77134
rect 586302 50218 586538 50454
rect 586622 50218 586858 50454
rect 586302 49898 586538 50134
rect 586622 49898 586858 50134
rect 586302 23218 586538 23454
rect 586622 23218 586858 23454
rect 586302 22898 586538 23134
rect 586622 22898 586858 23134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 701829 592650 701861
rect -8726 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 592650 701829
rect -8726 701509 592650 701593
rect -8726 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 592650 701509
rect -8726 701241 592650 701273
rect -8726 698454 592650 698486
rect -8726 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 592650 698454
rect -8726 698134 592650 698218
rect -8726 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 592650 698134
rect -8726 697866 592650 697898
rect -8726 674829 592650 674861
rect -8726 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 19952 674829
rect 20188 674593 25882 674829
rect 26118 674593 31813 674829
rect 32049 674593 47952 674829
rect 48188 674593 53882 674829
rect 54118 674593 59813 674829
rect 60049 674593 75952 674829
rect 76188 674593 81882 674829
rect 82118 674593 87813 674829
rect 88049 674593 103952 674829
rect 104188 674593 109882 674829
rect 110118 674593 115813 674829
rect 116049 674593 131952 674829
rect 132188 674593 137882 674829
rect 138118 674593 143813 674829
rect 144049 674593 159952 674829
rect 160188 674593 165882 674829
rect 166118 674593 171813 674829
rect 172049 674593 187952 674829
rect 188188 674593 193882 674829
rect 194118 674593 199813 674829
rect 200049 674593 215952 674829
rect 216188 674593 221882 674829
rect 222118 674593 227813 674829
rect 228049 674593 243952 674829
rect 244188 674593 249882 674829
rect 250118 674593 255813 674829
rect 256049 674593 271952 674829
rect 272188 674593 277882 674829
rect 278118 674593 283813 674829
rect 284049 674593 299952 674829
rect 300188 674593 305882 674829
rect 306118 674593 311813 674829
rect 312049 674593 327952 674829
rect 328188 674593 333882 674829
rect 334118 674593 339813 674829
rect 340049 674593 355952 674829
rect 356188 674593 361882 674829
rect 362118 674593 367813 674829
rect 368049 674593 383952 674829
rect 384188 674593 389882 674829
rect 390118 674593 395813 674829
rect 396049 674593 411952 674829
rect 412188 674593 417882 674829
rect 418118 674593 423813 674829
rect 424049 674593 439952 674829
rect 440188 674593 445882 674829
rect 446118 674593 451813 674829
rect 452049 674593 467952 674829
rect 468188 674593 473882 674829
rect 474118 674593 479813 674829
rect 480049 674593 495952 674829
rect 496188 674593 501882 674829
rect 502118 674593 507813 674829
rect 508049 674593 523952 674829
rect 524188 674593 529882 674829
rect 530118 674593 535813 674829
rect 536049 674593 551952 674829
rect 552188 674593 557882 674829
rect 558118 674593 563813 674829
rect 564049 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 592650 674829
rect -8726 674509 592650 674593
rect -8726 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 19952 674509
rect 20188 674273 25882 674509
rect 26118 674273 31813 674509
rect 32049 674273 47952 674509
rect 48188 674273 53882 674509
rect 54118 674273 59813 674509
rect 60049 674273 75952 674509
rect 76188 674273 81882 674509
rect 82118 674273 87813 674509
rect 88049 674273 103952 674509
rect 104188 674273 109882 674509
rect 110118 674273 115813 674509
rect 116049 674273 131952 674509
rect 132188 674273 137882 674509
rect 138118 674273 143813 674509
rect 144049 674273 159952 674509
rect 160188 674273 165882 674509
rect 166118 674273 171813 674509
rect 172049 674273 187952 674509
rect 188188 674273 193882 674509
rect 194118 674273 199813 674509
rect 200049 674273 215952 674509
rect 216188 674273 221882 674509
rect 222118 674273 227813 674509
rect 228049 674273 243952 674509
rect 244188 674273 249882 674509
rect 250118 674273 255813 674509
rect 256049 674273 271952 674509
rect 272188 674273 277882 674509
rect 278118 674273 283813 674509
rect 284049 674273 299952 674509
rect 300188 674273 305882 674509
rect 306118 674273 311813 674509
rect 312049 674273 327952 674509
rect 328188 674273 333882 674509
rect 334118 674273 339813 674509
rect 340049 674273 355952 674509
rect 356188 674273 361882 674509
rect 362118 674273 367813 674509
rect 368049 674273 383952 674509
rect 384188 674273 389882 674509
rect 390118 674273 395813 674509
rect 396049 674273 411952 674509
rect 412188 674273 417882 674509
rect 418118 674273 423813 674509
rect 424049 674273 439952 674509
rect 440188 674273 445882 674509
rect 446118 674273 451813 674509
rect 452049 674273 467952 674509
rect 468188 674273 473882 674509
rect 474118 674273 479813 674509
rect 480049 674273 495952 674509
rect 496188 674273 501882 674509
rect 502118 674273 507813 674509
rect 508049 674273 523952 674509
rect 524188 674273 529882 674509
rect 530118 674273 535813 674509
rect 536049 674273 551952 674509
rect 552188 674273 557882 674509
rect 558118 674273 563813 674509
rect 564049 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 592650 674509
rect -8726 674241 592650 674273
rect -8726 671454 592650 671486
rect -8726 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 22916 671454
rect 23152 671218 28847 671454
rect 29083 671218 50916 671454
rect 51152 671218 56847 671454
rect 57083 671218 78916 671454
rect 79152 671218 84847 671454
rect 85083 671218 106916 671454
rect 107152 671218 112847 671454
rect 113083 671218 134916 671454
rect 135152 671218 140847 671454
rect 141083 671218 162916 671454
rect 163152 671218 168847 671454
rect 169083 671218 190916 671454
rect 191152 671218 196847 671454
rect 197083 671218 218916 671454
rect 219152 671218 224847 671454
rect 225083 671218 246916 671454
rect 247152 671218 252847 671454
rect 253083 671218 274916 671454
rect 275152 671218 280847 671454
rect 281083 671218 302916 671454
rect 303152 671218 308847 671454
rect 309083 671218 330916 671454
rect 331152 671218 336847 671454
rect 337083 671218 358916 671454
rect 359152 671218 364847 671454
rect 365083 671218 386916 671454
rect 387152 671218 392847 671454
rect 393083 671218 414916 671454
rect 415152 671218 420847 671454
rect 421083 671218 442916 671454
rect 443152 671218 448847 671454
rect 449083 671218 470916 671454
rect 471152 671218 476847 671454
rect 477083 671218 498916 671454
rect 499152 671218 504847 671454
rect 505083 671218 526916 671454
rect 527152 671218 532847 671454
rect 533083 671218 554916 671454
rect 555152 671218 560847 671454
rect 561083 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 592650 671454
rect -8726 671134 592650 671218
rect -8726 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 22916 671134
rect 23152 670898 28847 671134
rect 29083 670898 50916 671134
rect 51152 670898 56847 671134
rect 57083 670898 78916 671134
rect 79152 670898 84847 671134
rect 85083 670898 106916 671134
rect 107152 670898 112847 671134
rect 113083 670898 134916 671134
rect 135152 670898 140847 671134
rect 141083 670898 162916 671134
rect 163152 670898 168847 671134
rect 169083 670898 190916 671134
rect 191152 670898 196847 671134
rect 197083 670898 218916 671134
rect 219152 670898 224847 671134
rect 225083 670898 246916 671134
rect 247152 670898 252847 671134
rect 253083 670898 274916 671134
rect 275152 670898 280847 671134
rect 281083 670898 302916 671134
rect 303152 670898 308847 671134
rect 309083 670898 330916 671134
rect 331152 670898 336847 671134
rect 337083 670898 358916 671134
rect 359152 670898 364847 671134
rect 365083 670898 386916 671134
rect 387152 670898 392847 671134
rect 393083 670898 414916 671134
rect 415152 670898 420847 671134
rect 421083 670898 442916 671134
rect 443152 670898 448847 671134
rect 449083 670898 470916 671134
rect 471152 670898 476847 671134
rect 477083 670898 498916 671134
rect 499152 670898 504847 671134
rect 505083 670898 526916 671134
rect 527152 670898 532847 671134
rect 533083 670898 554916 671134
rect 555152 670898 560847 671134
rect 561083 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 592650 671134
rect -8726 670866 592650 670898
rect -8726 647829 592650 647861
rect -8726 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 19952 647829
rect 20188 647593 25882 647829
rect 26118 647593 31813 647829
rect 32049 647593 47952 647829
rect 48188 647593 53882 647829
rect 54118 647593 59813 647829
rect 60049 647593 75952 647829
rect 76188 647593 81882 647829
rect 82118 647593 87813 647829
rect 88049 647593 103952 647829
rect 104188 647593 109882 647829
rect 110118 647593 115813 647829
rect 116049 647593 131952 647829
rect 132188 647593 137882 647829
rect 138118 647593 143813 647829
rect 144049 647593 159952 647829
rect 160188 647593 165882 647829
rect 166118 647593 171813 647829
rect 172049 647593 187952 647829
rect 188188 647593 193882 647829
rect 194118 647593 199813 647829
rect 200049 647593 215952 647829
rect 216188 647593 221882 647829
rect 222118 647593 227813 647829
rect 228049 647593 243952 647829
rect 244188 647593 249882 647829
rect 250118 647593 255813 647829
rect 256049 647593 271952 647829
rect 272188 647593 277882 647829
rect 278118 647593 283813 647829
rect 284049 647593 299952 647829
rect 300188 647593 305882 647829
rect 306118 647593 311813 647829
rect 312049 647593 327952 647829
rect 328188 647593 333882 647829
rect 334118 647593 339813 647829
rect 340049 647593 355952 647829
rect 356188 647593 361882 647829
rect 362118 647593 367813 647829
rect 368049 647593 383952 647829
rect 384188 647593 389882 647829
rect 390118 647593 395813 647829
rect 396049 647593 411952 647829
rect 412188 647593 417882 647829
rect 418118 647593 423813 647829
rect 424049 647593 439952 647829
rect 440188 647593 445882 647829
rect 446118 647593 451813 647829
rect 452049 647593 467952 647829
rect 468188 647593 473882 647829
rect 474118 647593 479813 647829
rect 480049 647593 495952 647829
rect 496188 647593 501882 647829
rect 502118 647593 507813 647829
rect 508049 647593 523952 647829
rect 524188 647593 529882 647829
rect 530118 647593 535813 647829
rect 536049 647593 551952 647829
rect 552188 647593 557882 647829
rect 558118 647593 563813 647829
rect 564049 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 592650 647829
rect -8726 647509 592650 647593
rect -8726 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 19952 647509
rect 20188 647273 25882 647509
rect 26118 647273 31813 647509
rect 32049 647273 47952 647509
rect 48188 647273 53882 647509
rect 54118 647273 59813 647509
rect 60049 647273 75952 647509
rect 76188 647273 81882 647509
rect 82118 647273 87813 647509
rect 88049 647273 103952 647509
rect 104188 647273 109882 647509
rect 110118 647273 115813 647509
rect 116049 647273 131952 647509
rect 132188 647273 137882 647509
rect 138118 647273 143813 647509
rect 144049 647273 159952 647509
rect 160188 647273 165882 647509
rect 166118 647273 171813 647509
rect 172049 647273 187952 647509
rect 188188 647273 193882 647509
rect 194118 647273 199813 647509
rect 200049 647273 215952 647509
rect 216188 647273 221882 647509
rect 222118 647273 227813 647509
rect 228049 647273 243952 647509
rect 244188 647273 249882 647509
rect 250118 647273 255813 647509
rect 256049 647273 271952 647509
rect 272188 647273 277882 647509
rect 278118 647273 283813 647509
rect 284049 647273 299952 647509
rect 300188 647273 305882 647509
rect 306118 647273 311813 647509
rect 312049 647273 327952 647509
rect 328188 647273 333882 647509
rect 334118 647273 339813 647509
rect 340049 647273 355952 647509
rect 356188 647273 361882 647509
rect 362118 647273 367813 647509
rect 368049 647273 383952 647509
rect 384188 647273 389882 647509
rect 390118 647273 395813 647509
rect 396049 647273 411952 647509
rect 412188 647273 417882 647509
rect 418118 647273 423813 647509
rect 424049 647273 439952 647509
rect 440188 647273 445882 647509
rect 446118 647273 451813 647509
rect 452049 647273 467952 647509
rect 468188 647273 473882 647509
rect 474118 647273 479813 647509
rect 480049 647273 495952 647509
rect 496188 647273 501882 647509
rect 502118 647273 507813 647509
rect 508049 647273 523952 647509
rect 524188 647273 529882 647509
rect 530118 647273 535813 647509
rect 536049 647273 551952 647509
rect 552188 647273 557882 647509
rect 558118 647273 563813 647509
rect 564049 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 592650 647509
rect -8726 647241 592650 647273
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 22916 644454
rect 23152 644218 28847 644454
rect 29083 644218 50916 644454
rect 51152 644218 56847 644454
rect 57083 644218 78916 644454
rect 79152 644218 84847 644454
rect 85083 644218 106916 644454
rect 107152 644218 112847 644454
rect 113083 644218 134916 644454
rect 135152 644218 140847 644454
rect 141083 644218 162916 644454
rect 163152 644218 168847 644454
rect 169083 644218 190916 644454
rect 191152 644218 196847 644454
rect 197083 644218 218916 644454
rect 219152 644218 224847 644454
rect 225083 644218 246916 644454
rect 247152 644218 252847 644454
rect 253083 644218 274916 644454
rect 275152 644218 280847 644454
rect 281083 644218 302916 644454
rect 303152 644218 308847 644454
rect 309083 644218 330916 644454
rect 331152 644218 336847 644454
rect 337083 644218 358916 644454
rect 359152 644218 364847 644454
rect 365083 644218 386916 644454
rect 387152 644218 392847 644454
rect 393083 644218 414916 644454
rect 415152 644218 420847 644454
rect 421083 644218 442916 644454
rect 443152 644218 448847 644454
rect 449083 644218 470916 644454
rect 471152 644218 476847 644454
rect 477083 644218 498916 644454
rect 499152 644218 504847 644454
rect 505083 644218 526916 644454
rect 527152 644218 532847 644454
rect 533083 644218 554916 644454
rect 555152 644218 560847 644454
rect 561083 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 22916 644134
rect 23152 643898 28847 644134
rect 29083 643898 50916 644134
rect 51152 643898 56847 644134
rect 57083 643898 78916 644134
rect 79152 643898 84847 644134
rect 85083 643898 106916 644134
rect 107152 643898 112847 644134
rect 113083 643898 134916 644134
rect 135152 643898 140847 644134
rect 141083 643898 162916 644134
rect 163152 643898 168847 644134
rect 169083 643898 190916 644134
rect 191152 643898 196847 644134
rect 197083 643898 218916 644134
rect 219152 643898 224847 644134
rect 225083 643898 246916 644134
rect 247152 643898 252847 644134
rect 253083 643898 274916 644134
rect 275152 643898 280847 644134
rect 281083 643898 302916 644134
rect 303152 643898 308847 644134
rect 309083 643898 330916 644134
rect 331152 643898 336847 644134
rect 337083 643898 358916 644134
rect 359152 643898 364847 644134
rect 365083 643898 386916 644134
rect 387152 643898 392847 644134
rect 393083 643898 414916 644134
rect 415152 643898 420847 644134
rect 421083 643898 442916 644134
rect 443152 643898 448847 644134
rect 449083 643898 470916 644134
rect 471152 643898 476847 644134
rect 477083 643898 498916 644134
rect 499152 643898 504847 644134
rect 505083 643898 526916 644134
rect 527152 643898 532847 644134
rect 533083 643898 554916 644134
rect 555152 643898 560847 644134
rect 561083 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 620829 592650 620861
rect -8726 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 19952 620829
rect 20188 620593 25882 620829
rect 26118 620593 31813 620829
rect 32049 620593 47952 620829
rect 48188 620593 53882 620829
rect 54118 620593 59813 620829
rect 60049 620593 75952 620829
rect 76188 620593 81882 620829
rect 82118 620593 87813 620829
rect 88049 620593 103952 620829
rect 104188 620593 109882 620829
rect 110118 620593 115813 620829
rect 116049 620593 131952 620829
rect 132188 620593 137882 620829
rect 138118 620593 143813 620829
rect 144049 620593 159952 620829
rect 160188 620593 165882 620829
rect 166118 620593 171813 620829
rect 172049 620593 187952 620829
rect 188188 620593 193882 620829
rect 194118 620593 199813 620829
rect 200049 620593 215952 620829
rect 216188 620593 221882 620829
rect 222118 620593 227813 620829
rect 228049 620593 243952 620829
rect 244188 620593 249882 620829
rect 250118 620593 255813 620829
rect 256049 620593 271952 620829
rect 272188 620593 277882 620829
rect 278118 620593 283813 620829
rect 284049 620593 299952 620829
rect 300188 620593 305882 620829
rect 306118 620593 311813 620829
rect 312049 620593 327952 620829
rect 328188 620593 333882 620829
rect 334118 620593 339813 620829
rect 340049 620593 355952 620829
rect 356188 620593 361882 620829
rect 362118 620593 367813 620829
rect 368049 620593 383952 620829
rect 384188 620593 389882 620829
rect 390118 620593 395813 620829
rect 396049 620593 411952 620829
rect 412188 620593 417882 620829
rect 418118 620593 423813 620829
rect 424049 620593 439952 620829
rect 440188 620593 445882 620829
rect 446118 620593 451813 620829
rect 452049 620593 467952 620829
rect 468188 620593 473882 620829
rect 474118 620593 479813 620829
rect 480049 620593 495952 620829
rect 496188 620593 501882 620829
rect 502118 620593 507813 620829
rect 508049 620593 523952 620829
rect 524188 620593 529882 620829
rect 530118 620593 535813 620829
rect 536049 620593 551952 620829
rect 552188 620593 557882 620829
rect 558118 620593 563813 620829
rect 564049 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 592650 620829
rect -8726 620509 592650 620593
rect -8726 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 19952 620509
rect 20188 620273 25882 620509
rect 26118 620273 31813 620509
rect 32049 620273 47952 620509
rect 48188 620273 53882 620509
rect 54118 620273 59813 620509
rect 60049 620273 75952 620509
rect 76188 620273 81882 620509
rect 82118 620273 87813 620509
rect 88049 620273 103952 620509
rect 104188 620273 109882 620509
rect 110118 620273 115813 620509
rect 116049 620273 131952 620509
rect 132188 620273 137882 620509
rect 138118 620273 143813 620509
rect 144049 620273 159952 620509
rect 160188 620273 165882 620509
rect 166118 620273 171813 620509
rect 172049 620273 187952 620509
rect 188188 620273 193882 620509
rect 194118 620273 199813 620509
rect 200049 620273 215952 620509
rect 216188 620273 221882 620509
rect 222118 620273 227813 620509
rect 228049 620273 243952 620509
rect 244188 620273 249882 620509
rect 250118 620273 255813 620509
rect 256049 620273 271952 620509
rect 272188 620273 277882 620509
rect 278118 620273 283813 620509
rect 284049 620273 299952 620509
rect 300188 620273 305882 620509
rect 306118 620273 311813 620509
rect 312049 620273 327952 620509
rect 328188 620273 333882 620509
rect 334118 620273 339813 620509
rect 340049 620273 355952 620509
rect 356188 620273 361882 620509
rect 362118 620273 367813 620509
rect 368049 620273 383952 620509
rect 384188 620273 389882 620509
rect 390118 620273 395813 620509
rect 396049 620273 411952 620509
rect 412188 620273 417882 620509
rect 418118 620273 423813 620509
rect 424049 620273 439952 620509
rect 440188 620273 445882 620509
rect 446118 620273 451813 620509
rect 452049 620273 467952 620509
rect 468188 620273 473882 620509
rect 474118 620273 479813 620509
rect 480049 620273 495952 620509
rect 496188 620273 501882 620509
rect 502118 620273 507813 620509
rect 508049 620273 523952 620509
rect 524188 620273 529882 620509
rect 530118 620273 535813 620509
rect 536049 620273 551952 620509
rect 552188 620273 557882 620509
rect 558118 620273 563813 620509
rect 564049 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 592650 620509
rect -8726 620241 592650 620273
rect -8726 617454 592650 617486
rect -8726 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 22916 617454
rect 23152 617218 28847 617454
rect 29083 617218 50916 617454
rect 51152 617218 56847 617454
rect 57083 617218 78916 617454
rect 79152 617218 84847 617454
rect 85083 617218 106916 617454
rect 107152 617218 112847 617454
rect 113083 617218 134916 617454
rect 135152 617218 140847 617454
rect 141083 617218 162916 617454
rect 163152 617218 168847 617454
rect 169083 617218 190916 617454
rect 191152 617218 196847 617454
rect 197083 617218 218916 617454
rect 219152 617218 224847 617454
rect 225083 617218 246916 617454
rect 247152 617218 252847 617454
rect 253083 617218 274916 617454
rect 275152 617218 280847 617454
rect 281083 617218 302916 617454
rect 303152 617218 308847 617454
rect 309083 617218 330916 617454
rect 331152 617218 336847 617454
rect 337083 617218 358916 617454
rect 359152 617218 364847 617454
rect 365083 617218 386916 617454
rect 387152 617218 392847 617454
rect 393083 617218 414916 617454
rect 415152 617218 420847 617454
rect 421083 617218 442916 617454
rect 443152 617218 448847 617454
rect 449083 617218 470916 617454
rect 471152 617218 476847 617454
rect 477083 617218 498916 617454
rect 499152 617218 504847 617454
rect 505083 617218 526916 617454
rect 527152 617218 532847 617454
rect 533083 617218 554916 617454
rect 555152 617218 560847 617454
rect 561083 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 592650 617454
rect -8726 617134 592650 617218
rect -8726 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 22916 617134
rect 23152 616898 28847 617134
rect 29083 616898 50916 617134
rect 51152 616898 56847 617134
rect 57083 616898 78916 617134
rect 79152 616898 84847 617134
rect 85083 616898 106916 617134
rect 107152 616898 112847 617134
rect 113083 616898 134916 617134
rect 135152 616898 140847 617134
rect 141083 616898 162916 617134
rect 163152 616898 168847 617134
rect 169083 616898 190916 617134
rect 191152 616898 196847 617134
rect 197083 616898 218916 617134
rect 219152 616898 224847 617134
rect 225083 616898 246916 617134
rect 247152 616898 252847 617134
rect 253083 616898 274916 617134
rect 275152 616898 280847 617134
rect 281083 616898 302916 617134
rect 303152 616898 308847 617134
rect 309083 616898 330916 617134
rect 331152 616898 336847 617134
rect 337083 616898 358916 617134
rect 359152 616898 364847 617134
rect 365083 616898 386916 617134
rect 387152 616898 392847 617134
rect 393083 616898 414916 617134
rect 415152 616898 420847 617134
rect 421083 616898 442916 617134
rect 443152 616898 448847 617134
rect 449083 616898 470916 617134
rect 471152 616898 476847 617134
rect 477083 616898 498916 617134
rect 499152 616898 504847 617134
rect 505083 616898 526916 617134
rect 527152 616898 532847 617134
rect 533083 616898 554916 617134
rect 555152 616898 560847 617134
rect 561083 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 592650 617134
rect -8726 616866 592650 616898
rect -8726 593829 592650 593861
rect -8726 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 19952 593829
rect 20188 593593 25882 593829
rect 26118 593593 31813 593829
rect 32049 593593 47952 593829
rect 48188 593593 53882 593829
rect 54118 593593 59813 593829
rect 60049 593593 75952 593829
rect 76188 593593 81882 593829
rect 82118 593593 87813 593829
rect 88049 593593 103952 593829
rect 104188 593593 109882 593829
rect 110118 593593 115813 593829
rect 116049 593593 131952 593829
rect 132188 593593 137882 593829
rect 138118 593593 143813 593829
rect 144049 593593 159952 593829
rect 160188 593593 165882 593829
rect 166118 593593 171813 593829
rect 172049 593593 187952 593829
rect 188188 593593 193882 593829
rect 194118 593593 199813 593829
rect 200049 593593 215952 593829
rect 216188 593593 221882 593829
rect 222118 593593 227813 593829
rect 228049 593593 243952 593829
rect 244188 593593 249882 593829
rect 250118 593593 255813 593829
rect 256049 593593 271952 593829
rect 272188 593593 277882 593829
rect 278118 593593 283813 593829
rect 284049 593593 299952 593829
rect 300188 593593 305882 593829
rect 306118 593593 311813 593829
rect 312049 593593 327952 593829
rect 328188 593593 333882 593829
rect 334118 593593 339813 593829
rect 340049 593593 355952 593829
rect 356188 593593 361882 593829
rect 362118 593593 367813 593829
rect 368049 593593 383952 593829
rect 384188 593593 389882 593829
rect 390118 593593 395813 593829
rect 396049 593593 411952 593829
rect 412188 593593 417882 593829
rect 418118 593593 423813 593829
rect 424049 593593 439952 593829
rect 440188 593593 445882 593829
rect 446118 593593 451813 593829
rect 452049 593593 467952 593829
rect 468188 593593 473882 593829
rect 474118 593593 479813 593829
rect 480049 593593 495952 593829
rect 496188 593593 501882 593829
rect 502118 593593 507813 593829
rect 508049 593593 523952 593829
rect 524188 593593 529882 593829
rect 530118 593593 535813 593829
rect 536049 593593 551952 593829
rect 552188 593593 557882 593829
rect 558118 593593 563813 593829
rect 564049 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 592650 593829
rect -8726 593509 592650 593593
rect -8726 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 19952 593509
rect 20188 593273 25882 593509
rect 26118 593273 31813 593509
rect 32049 593273 47952 593509
rect 48188 593273 53882 593509
rect 54118 593273 59813 593509
rect 60049 593273 75952 593509
rect 76188 593273 81882 593509
rect 82118 593273 87813 593509
rect 88049 593273 103952 593509
rect 104188 593273 109882 593509
rect 110118 593273 115813 593509
rect 116049 593273 131952 593509
rect 132188 593273 137882 593509
rect 138118 593273 143813 593509
rect 144049 593273 159952 593509
rect 160188 593273 165882 593509
rect 166118 593273 171813 593509
rect 172049 593273 187952 593509
rect 188188 593273 193882 593509
rect 194118 593273 199813 593509
rect 200049 593273 215952 593509
rect 216188 593273 221882 593509
rect 222118 593273 227813 593509
rect 228049 593273 243952 593509
rect 244188 593273 249882 593509
rect 250118 593273 255813 593509
rect 256049 593273 271952 593509
rect 272188 593273 277882 593509
rect 278118 593273 283813 593509
rect 284049 593273 299952 593509
rect 300188 593273 305882 593509
rect 306118 593273 311813 593509
rect 312049 593273 327952 593509
rect 328188 593273 333882 593509
rect 334118 593273 339813 593509
rect 340049 593273 355952 593509
rect 356188 593273 361882 593509
rect 362118 593273 367813 593509
rect 368049 593273 383952 593509
rect 384188 593273 389882 593509
rect 390118 593273 395813 593509
rect 396049 593273 411952 593509
rect 412188 593273 417882 593509
rect 418118 593273 423813 593509
rect 424049 593273 439952 593509
rect 440188 593273 445882 593509
rect 446118 593273 451813 593509
rect 452049 593273 467952 593509
rect 468188 593273 473882 593509
rect 474118 593273 479813 593509
rect 480049 593273 495952 593509
rect 496188 593273 501882 593509
rect 502118 593273 507813 593509
rect 508049 593273 523952 593509
rect 524188 593273 529882 593509
rect 530118 593273 535813 593509
rect 536049 593273 551952 593509
rect 552188 593273 557882 593509
rect 558118 593273 563813 593509
rect 564049 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 592650 593509
rect -8726 593241 592650 593273
rect -8726 590454 592650 590486
rect -8726 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 22916 590454
rect 23152 590218 28847 590454
rect 29083 590218 50916 590454
rect 51152 590218 56847 590454
rect 57083 590218 78916 590454
rect 79152 590218 84847 590454
rect 85083 590218 106916 590454
rect 107152 590218 112847 590454
rect 113083 590218 134916 590454
rect 135152 590218 140847 590454
rect 141083 590218 162916 590454
rect 163152 590218 168847 590454
rect 169083 590218 190916 590454
rect 191152 590218 196847 590454
rect 197083 590218 218916 590454
rect 219152 590218 224847 590454
rect 225083 590218 246916 590454
rect 247152 590218 252847 590454
rect 253083 590218 274916 590454
rect 275152 590218 280847 590454
rect 281083 590218 302916 590454
rect 303152 590218 308847 590454
rect 309083 590218 330916 590454
rect 331152 590218 336847 590454
rect 337083 590218 358916 590454
rect 359152 590218 364847 590454
rect 365083 590218 386916 590454
rect 387152 590218 392847 590454
rect 393083 590218 414916 590454
rect 415152 590218 420847 590454
rect 421083 590218 442916 590454
rect 443152 590218 448847 590454
rect 449083 590218 470916 590454
rect 471152 590218 476847 590454
rect 477083 590218 498916 590454
rect 499152 590218 504847 590454
rect 505083 590218 526916 590454
rect 527152 590218 532847 590454
rect 533083 590218 554916 590454
rect 555152 590218 560847 590454
rect 561083 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 592650 590454
rect -8726 590134 592650 590218
rect -8726 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 22916 590134
rect 23152 589898 28847 590134
rect 29083 589898 50916 590134
rect 51152 589898 56847 590134
rect 57083 589898 78916 590134
rect 79152 589898 84847 590134
rect 85083 589898 106916 590134
rect 107152 589898 112847 590134
rect 113083 589898 134916 590134
rect 135152 589898 140847 590134
rect 141083 589898 162916 590134
rect 163152 589898 168847 590134
rect 169083 589898 190916 590134
rect 191152 589898 196847 590134
rect 197083 589898 218916 590134
rect 219152 589898 224847 590134
rect 225083 589898 246916 590134
rect 247152 589898 252847 590134
rect 253083 589898 274916 590134
rect 275152 589898 280847 590134
rect 281083 589898 302916 590134
rect 303152 589898 308847 590134
rect 309083 589898 330916 590134
rect 331152 589898 336847 590134
rect 337083 589898 358916 590134
rect 359152 589898 364847 590134
rect 365083 589898 386916 590134
rect 387152 589898 392847 590134
rect 393083 589898 414916 590134
rect 415152 589898 420847 590134
rect 421083 589898 442916 590134
rect 443152 589898 448847 590134
rect 449083 589898 470916 590134
rect 471152 589898 476847 590134
rect 477083 589898 498916 590134
rect 499152 589898 504847 590134
rect 505083 589898 526916 590134
rect 527152 589898 532847 590134
rect 533083 589898 554916 590134
rect 555152 589898 560847 590134
rect 561083 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 592650 590134
rect -8726 589866 592650 589898
rect -8726 566829 592650 566861
rect -8726 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 19952 566829
rect 20188 566593 25882 566829
rect 26118 566593 31813 566829
rect 32049 566593 47952 566829
rect 48188 566593 53882 566829
rect 54118 566593 59813 566829
rect 60049 566593 75952 566829
rect 76188 566593 81882 566829
rect 82118 566593 87813 566829
rect 88049 566593 103952 566829
rect 104188 566593 109882 566829
rect 110118 566593 115813 566829
rect 116049 566593 131952 566829
rect 132188 566593 137882 566829
rect 138118 566593 143813 566829
rect 144049 566593 159952 566829
rect 160188 566593 165882 566829
rect 166118 566593 171813 566829
rect 172049 566593 187952 566829
rect 188188 566593 193882 566829
rect 194118 566593 199813 566829
rect 200049 566593 215952 566829
rect 216188 566593 221882 566829
rect 222118 566593 227813 566829
rect 228049 566593 243952 566829
rect 244188 566593 249882 566829
rect 250118 566593 255813 566829
rect 256049 566593 271952 566829
rect 272188 566593 277882 566829
rect 278118 566593 283813 566829
rect 284049 566593 299952 566829
rect 300188 566593 305882 566829
rect 306118 566593 311813 566829
rect 312049 566593 327952 566829
rect 328188 566593 333882 566829
rect 334118 566593 339813 566829
rect 340049 566593 355952 566829
rect 356188 566593 361882 566829
rect 362118 566593 367813 566829
rect 368049 566593 383952 566829
rect 384188 566593 389882 566829
rect 390118 566593 395813 566829
rect 396049 566593 411952 566829
rect 412188 566593 417882 566829
rect 418118 566593 423813 566829
rect 424049 566593 439952 566829
rect 440188 566593 445882 566829
rect 446118 566593 451813 566829
rect 452049 566593 467952 566829
rect 468188 566593 473882 566829
rect 474118 566593 479813 566829
rect 480049 566593 495952 566829
rect 496188 566593 501882 566829
rect 502118 566593 507813 566829
rect 508049 566593 523952 566829
rect 524188 566593 529882 566829
rect 530118 566593 535813 566829
rect 536049 566593 551952 566829
rect 552188 566593 557882 566829
rect 558118 566593 563813 566829
rect 564049 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 592650 566829
rect -8726 566509 592650 566593
rect -8726 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 19952 566509
rect 20188 566273 25882 566509
rect 26118 566273 31813 566509
rect 32049 566273 47952 566509
rect 48188 566273 53882 566509
rect 54118 566273 59813 566509
rect 60049 566273 75952 566509
rect 76188 566273 81882 566509
rect 82118 566273 87813 566509
rect 88049 566273 103952 566509
rect 104188 566273 109882 566509
rect 110118 566273 115813 566509
rect 116049 566273 131952 566509
rect 132188 566273 137882 566509
rect 138118 566273 143813 566509
rect 144049 566273 159952 566509
rect 160188 566273 165882 566509
rect 166118 566273 171813 566509
rect 172049 566273 187952 566509
rect 188188 566273 193882 566509
rect 194118 566273 199813 566509
rect 200049 566273 215952 566509
rect 216188 566273 221882 566509
rect 222118 566273 227813 566509
rect 228049 566273 243952 566509
rect 244188 566273 249882 566509
rect 250118 566273 255813 566509
rect 256049 566273 271952 566509
rect 272188 566273 277882 566509
rect 278118 566273 283813 566509
rect 284049 566273 299952 566509
rect 300188 566273 305882 566509
rect 306118 566273 311813 566509
rect 312049 566273 327952 566509
rect 328188 566273 333882 566509
rect 334118 566273 339813 566509
rect 340049 566273 355952 566509
rect 356188 566273 361882 566509
rect 362118 566273 367813 566509
rect 368049 566273 383952 566509
rect 384188 566273 389882 566509
rect 390118 566273 395813 566509
rect 396049 566273 411952 566509
rect 412188 566273 417882 566509
rect 418118 566273 423813 566509
rect 424049 566273 439952 566509
rect 440188 566273 445882 566509
rect 446118 566273 451813 566509
rect 452049 566273 467952 566509
rect 468188 566273 473882 566509
rect 474118 566273 479813 566509
rect 480049 566273 495952 566509
rect 496188 566273 501882 566509
rect 502118 566273 507813 566509
rect 508049 566273 523952 566509
rect 524188 566273 529882 566509
rect 530118 566273 535813 566509
rect 536049 566273 551952 566509
rect 552188 566273 557882 566509
rect 558118 566273 563813 566509
rect 564049 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 592650 566509
rect -8726 566241 592650 566273
rect -8726 563454 592650 563486
rect -8726 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 22916 563454
rect 23152 563218 28847 563454
rect 29083 563218 50916 563454
rect 51152 563218 56847 563454
rect 57083 563218 78916 563454
rect 79152 563218 84847 563454
rect 85083 563218 106916 563454
rect 107152 563218 112847 563454
rect 113083 563218 134916 563454
rect 135152 563218 140847 563454
rect 141083 563218 162916 563454
rect 163152 563218 168847 563454
rect 169083 563218 190916 563454
rect 191152 563218 196847 563454
rect 197083 563218 218916 563454
rect 219152 563218 224847 563454
rect 225083 563218 246916 563454
rect 247152 563218 252847 563454
rect 253083 563218 274916 563454
rect 275152 563218 280847 563454
rect 281083 563218 302916 563454
rect 303152 563218 308847 563454
rect 309083 563218 330916 563454
rect 331152 563218 336847 563454
rect 337083 563218 358916 563454
rect 359152 563218 364847 563454
rect 365083 563218 386916 563454
rect 387152 563218 392847 563454
rect 393083 563218 414916 563454
rect 415152 563218 420847 563454
rect 421083 563218 442916 563454
rect 443152 563218 448847 563454
rect 449083 563218 470916 563454
rect 471152 563218 476847 563454
rect 477083 563218 498916 563454
rect 499152 563218 504847 563454
rect 505083 563218 526916 563454
rect 527152 563218 532847 563454
rect 533083 563218 554916 563454
rect 555152 563218 560847 563454
rect 561083 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 592650 563454
rect -8726 563134 592650 563218
rect -8726 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 22916 563134
rect 23152 562898 28847 563134
rect 29083 562898 50916 563134
rect 51152 562898 56847 563134
rect 57083 562898 78916 563134
rect 79152 562898 84847 563134
rect 85083 562898 106916 563134
rect 107152 562898 112847 563134
rect 113083 562898 134916 563134
rect 135152 562898 140847 563134
rect 141083 562898 162916 563134
rect 163152 562898 168847 563134
rect 169083 562898 190916 563134
rect 191152 562898 196847 563134
rect 197083 562898 218916 563134
rect 219152 562898 224847 563134
rect 225083 562898 246916 563134
rect 247152 562898 252847 563134
rect 253083 562898 274916 563134
rect 275152 562898 280847 563134
rect 281083 562898 302916 563134
rect 303152 562898 308847 563134
rect 309083 562898 330916 563134
rect 331152 562898 336847 563134
rect 337083 562898 358916 563134
rect 359152 562898 364847 563134
rect 365083 562898 386916 563134
rect 387152 562898 392847 563134
rect 393083 562898 414916 563134
rect 415152 562898 420847 563134
rect 421083 562898 442916 563134
rect 443152 562898 448847 563134
rect 449083 562898 470916 563134
rect 471152 562898 476847 563134
rect 477083 562898 498916 563134
rect 499152 562898 504847 563134
rect 505083 562898 526916 563134
rect 527152 562898 532847 563134
rect 533083 562898 554916 563134
rect 555152 562898 560847 563134
rect 561083 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 592650 563134
rect -8726 562866 592650 562898
rect -8726 539829 592650 539861
rect -8726 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 19952 539829
rect 20188 539593 25882 539829
rect 26118 539593 31813 539829
rect 32049 539593 47952 539829
rect 48188 539593 53882 539829
rect 54118 539593 59813 539829
rect 60049 539593 75952 539829
rect 76188 539593 81882 539829
rect 82118 539593 87813 539829
rect 88049 539593 103952 539829
rect 104188 539593 109882 539829
rect 110118 539593 115813 539829
rect 116049 539593 131952 539829
rect 132188 539593 137882 539829
rect 138118 539593 143813 539829
rect 144049 539593 159952 539829
rect 160188 539593 165882 539829
rect 166118 539593 171813 539829
rect 172049 539593 187952 539829
rect 188188 539593 193882 539829
rect 194118 539593 199813 539829
rect 200049 539593 215952 539829
rect 216188 539593 221882 539829
rect 222118 539593 227813 539829
rect 228049 539593 243952 539829
rect 244188 539593 249882 539829
rect 250118 539593 255813 539829
rect 256049 539593 271952 539829
rect 272188 539593 277882 539829
rect 278118 539593 283813 539829
rect 284049 539593 299952 539829
rect 300188 539593 305882 539829
rect 306118 539593 311813 539829
rect 312049 539593 327952 539829
rect 328188 539593 333882 539829
rect 334118 539593 339813 539829
rect 340049 539593 355952 539829
rect 356188 539593 361882 539829
rect 362118 539593 367813 539829
rect 368049 539593 383952 539829
rect 384188 539593 389882 539829
rect 390118 539593 395813 539829
rect 396049 539593 411952 539829
rect 412188 539593 417882 539829
rect 418118 539593 423813 539829
rect 424049 539593 439952 539829
rect 440188 539593 445882 539829
rect 446118 539593 451813 539829
rect 452049 539593 467952 539829
rect 468188 539593 473882 539829
rect 474118 539593 479813 539829
rect 480049 539593 495952 539829
rect 496188 539593 501882 539829
rect 502118 539593 507813 539829
rect 508049 539593 523952 539829
rect 524188 539593 529882 539829
rect 530118 539593 535813 539829
rect 536049 539593 551952 539829
rect 552188 539593 557882 539829
rect 558118 539593 563813 539829
rect 564049 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 592650 539829
rect -8726 539509 592650 539593
rect -8726 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 19952 539509
rect 20188 539273 25882 539509
rect 26118 539273 31813 539509
rect 32049 539273 47952 539509
rect 48188 539273 53882 539509
rect 54118 539273 59813 539509
rect 60049 539273 75952 539509
rect 76188 539273 81882 539509
rect 82118 539273 87813 539509
rect 88049 539273 103952 539509
rect 104188 539273 109882 539509
rect 110118 539273 115813 539509
rect 116049 539273 131952 539509
rect 132188 539273 137882 539509
rect 138118 539273 143813 539509
rect 144049 539273 159952 539509
rect 160188 539273 165882 539509
rect 166118 539273 171813 539509
rect 172049 539273 187952 539509
rect 188188 539273 193882 539509
rect 194118 539273 199813 539509
rect 200049 539273 215952 539509
rect 216188 539273 221882 539509
rect 222118 539273 227813 539509
rect 228049 539273 243952 539509
rect 244188 539273 249882 539509
rect 250118 539273 255813 539509
rect 256049 539273 271952 539509
rect 272188 539273 277882 539509
rect 278118 539273 283813 539509
rect 284049 539273 299952 539509
rect 300188 539273 305882 539509
rect 306118 539273 311813 539509
rect 312049 539273 327952 539509
rect 328188 539273 333882 539509
rect 334118 539273 339813 539509
rect 340049 539273 355952 539509
rect 356188 539273 361882 539509
rect 362118 539273 367813 539509
rect 368049 539273 383952 539509
rect 384188 539273 389882 539509
rect 390118 539273 395813 539509
rect 396049 539273 411952 539509
rect 412188 539273 417882 539509
rect 418118 539273 423813 539509
rect 424049 539273 439952 539509
rect 440188 539273 445882 539509
rect 446118 539273 451813 539509
rect 452049 539273 467952 539509
rect 468188 539273 473882 539509
rect 474118 539273 479813 539509
rect 480049 539273 495952 539509
rect 496188 539273 501882 539509
rect 502118 539273 507813 539509
rect 508049 539273 523952 539509
rect 524188 539273 529882 539509
rect 530118 539273 535813 539509
rect 536049 539273 551952 539509
rect 552188 539273 557882 539509
rect 558118 539273 563813 539509
rect 564049 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 592650 539509
rect -8726 539241 592650 539273
rect -8726 536454 592650 536486
rect -8726 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 22916 536454
rect 23152 536218 28847 536454
rect 29083 536218 50916 536454
rect 51152 536218 56847 536454
rect 57083 536218 78916 536454
rect 79152 536218 84847 536454
rect 85083 536218 106916 536454
rect 107152 536218 112847 536454
rect 113083 536218 134916 536454
rect 135152 536218 140847 536454
rect 141083 536218 162916 536454
rect 163152 536218 168847 536454
rect 169083 536218 190916 536454
rect 191152 536218 196847 536454
rect 197083 536218 218916 536454
rect 219152 536218 224847 536454
rect 225083 536218 246916 536454
rect 247152 536218 252847 536454
rect 253083 536218 274916 536454
rect 275152 536218 280847 536454
rect 281083 536218 302916 536454
rect 303152 536218 308847 536454
rect 309083 536218 330916 536454
rect 331152 536218 336847 536454
rect 337083 536218 358916 536454
rect 359152 536218 364847 536454
rect 365083 536218 386916 536454
rect 387152 536218 392847 536454
rect 393083 536218 414916 536454
rect 415152 536218 420847 536454
rect 421083 536218 442916 536454
rect 443152 536218 448847 536454
rect 449083 536218 470916 536454
rect 471152 536218 476847 536454
rect 477083 536218 498916 536454
rect 499152 536218 504847 536454
rect 505083 536218 526916 536454
rect 527152 536218 532847 536454
rect 533083 536218 554916 536454
rect 555152 536218 560847 536454
rect 561083 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 592650 536454
rect -8726 536134 592650 536218
rect -8726 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 22916 536134
rect 23152 535898 28847 536134
rect 29083 535898 50916 536134
rect 51152 535898 56847 536134
rect 57083 535898 78916 536134
rect 79152 535898 84847 536134
rect 85083 535898 106916 536134
rect 107152 535898 112847 536134
rect 113083 535898 134916 536134
rect 135152 535898 140847 536134
rect 141083 535898 162916 536134
rect 163152 535898 168847 536134
rect 169083 535898 190916 536134
rect 191152 535898 196847 536134
rect 197083 535898 218916 536134
rect 219152 535898 224847 536134
rect 225083 535898 246916 536134
rect 247152 535898 252847 536134
rect 253083 535898 274916 536134
rect 275152 535898 280847 536134
rect 281083 535898 302916 536134
rect 303152 535898 308847 536134
rect 309083 535898 330916 536134
rect 331152 535898 336847 536134
rect 337083 535898 358916 536134
rect 359152 535898 364847 536134
rect 365083 535898 386916 536134
rect 387152 535898 392847 536134
rect 393083 535898 414916 536134
rect 415152 535898 420847 536134
rect 421083 535898 442916 536134
rect 443152 535898 448847 536134
rect 449083 535898 470916 536134
rect 471152 535898 476847 536134
rect 477083 535898 498916 536134
rect 499152 535898 504847 536134
rect 505083 535898 526916 536134
rect 527152 535898 532847 536134
rect 533083 535898 554916 536134
rect 555152 535898 560847 536134
rect 561083 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 592650 536134
rect -8726 535866 592650 535898
rect -8726 512829 592650 512861
rect -8726 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 19952 512829
rect 20188 512593 25882 512829
rect 26118 512593 31813 512829
rect 32049 512593 47952 512829
rect 48188 512593 53882 512829
rect 54118 512593 59813 512829
rect 60049 512593 75952 512829
rect 76188 512593 81882 512829
rect 82118 512593 87813 512829
rect 88049 512593 103952 512829
rect 104188 512593 109882 512829
rect 110118 512593 115813 512829
rect 116049 512593 131952 512829
rect 132188 512593 137882 512829
rect 138118 512593 143813 512829
rect 144049 512593 159952 512829
rect 160188 512593 165882 512829
rect 166118 512593 171813 512829
rect 172049 512593 187952 512829
rect 188188 512593 193882 512829
rect 194118 512593 199813 512829
rect 200049 512593 215952 512829
rect 216188 512593 221882 512829
rect 222118 512593 227813 512829
rect 228049 512593 243952 512829
rect 244188 512593 249882 512829
rect 250118 512593 255813 512829
rect 256049 512593 271952 512829
rect 272188 512593 277882 512829
rect 278118 512593 283813 512829
rect 284049 512593 299952 512829
rect 300188 512593 305882 512829
rect 306118 512593 311813 512829
rect 312049 512593 327952 512829
rect 328188 512593 333882 512829
rect 334118 512593 339813 512829
rect 340049 512593 355952 512829
rect 356188 512593 361882 512829
rect 362118 512593 367813 512829
rect 368049 512593 383952 512829
rect 384188 512593 389882 512829
rect 390118 512593 395813 512829
rect 396049 512593 411952 512829
rect 412188 512593 417882 512829
rect 418118 512593 423813 512829
rect 424049 512593 439952 512829
rect 440188 512593 445882 512829
rect 446118 512593 451813 512829
rect 452049 512593 467952 512829
rect 468188 512593 473882 512829
rect 474118 512593 479813 512829
rect 480049 512593 495952 512829
rect 496188 512593 501882 512829
rect 502118 512593 507813 512829
rect 508049 512593 523952 512829
rect 524188 512593 529882 512829
rect 530118 512593 535813 512829
rect 536049 512593 551952 512829
rect 552188 512593 557882 512829
rect 558118 512593 563813 512829
rect 564049 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 592650 512829
rect -8726 512509 592650 512593
rect -8726 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 19952 512509
rect 20188 512273 25882 512509
rect 26118 512273 31813 512509
rect 32049 512273 47952 512509
rect 48188 512273 53882 512509
rect 54118 512273 59813 512509
rect 60049 512273 75952 512509
rect 76188 512273 81882 512509
rect 82118 512273 87813 512509
rect 88049 512273 103952 512509
rect 104188 512273 109882 512509
rect 110118 512273 115813 512509
rect 116049 512273 131952 512509
rect 132188 512273 137882 512509
rect 138118 512273 143813 512509
rect 144049 512273 159952 512509
rect 160188 512273 165882 512509
rect 166118 512273 171813 512509
rect 172049 512273 187952 512509
rect 188188 512273 193882 512509
rect 194118 512273 199813 512509
rect 200049 512273 215952 512509
rect 216188 512273 221882 512509
rect 222118 512273 227813 512509
rect 228049 512273 243952 512509
rect 244188 512273 249882 512509
rect 250118 512273 255813 512509
rect 256049 512273 271952 512509
rect 272188 512273 277882 512509
rect 278118 512273 283813 512509
rect 284049 512273 299952 512509
rect 300188 512273 305882 512509
rect 306118 512273 311813 512509
rect 312049 512273 327952 512509
rect 328188 512273 333882 512509
rect 334118 512273 339813 512509
rect 340049 512273 355952 512509
rect 356188 512273 361882 512509
rect 362118 512273 367813 512509
rect 368049 512273 383952 512509
rect 384188 512273 389882 512509
rect 390118 512273 395813 512509
rect 396049 512273 411952 512509
rect 412188 512273 417882 512509
rect 418118 512273 423813 512509
rect 424049 512273 439952 512509
rect 440188 512273 445882 512509
rect 446118 512273 451813 512509
rect 452049 512273 467952 512509
rect 468188 512273 473882 512509
rect 474118 512273 479813 512509
rect 480049 512273 495952 512509
rect 496188 512273 501882 512509
rect 502118 512273 507813 512509
rect 508049 512273 523952 512509
rect 524188 512273 529882 512509
rect 530118 512273 535813 512509
rect 536049 512273 551952 512509
rect 552188 512273 557882 512509
rect 558118 512273 563813 512509
rect 564049 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 592650 512509
rect -8726 512241 592650 512273
rect -8726 509454 592650 509486
rect -8726 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 22916 509454
rect 23152 509218 28847 509454
rect 29083 509218 50916 509454
rect 51152 509218 56847 509454
rect 57083 509218 78916 509454
rect 79152 509218 84847 509454
rect 85083 509218 106916 509454
rect 107152 509218 112847 509454
rect 113083 509218 134916 509454
rect 135152 509218 140847 509454
rect 141083 509218 162916 509454
rect 163152 509218 168847 509454
rect 169083 509218 190916 509454
rect 191152 509218 196847 509454
rect 197083 509218 218916 509454
rect 219152 509218 224847 509454
rect 225083 509218 246916 509454
rect 247152 509218 252847 509454
rect 253083 509218 274916 509454
rect 275152 509218 280847 509454
rect 281083 509218 302916 509454
rect 303152 509218 308847 509454
rect 309083 509218 330916 509454
rect 331152 509218 336847 509454
rect 337083 509218 358916 509454
rect 359152 509218 364847 509454
rect 365083 509218 386916 509454
rect 387152 509218 392847 509454
rect 393083 509218 414916 509454
rect 415152 509218 420847 509454
rect 421083 509218 442916 509454
rect 443152 509218 448847 509454
rect 449083 509218 470916 509454
rect 471152 509218 476847 509454
rect 477083 509218 498916 509454
rect 499152 509218 504847 509454
rect 505083 509218 526916 509454
rect 527152 509218 532847 509454
rect 533083 509218 554916 509454
rect 555152 509218 560847 509454
rect 561083 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 592650 509454
rect -8726 509134 592650 509218
rect -8726 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 22916 509134
rect 23152 508898 28847 509134
rect 29083 508898 50916 509134
rect 51152 508898 56847 509134
rect 57083 508898 78916 509134
rect 79152 508898 84847 509134
rect 85083 508898 106916 509134
rect 107152 508898 112847 509134
rect 113083 508898 134916 509134
rect 135152 508898 140847 509134
rect 141083 508898 162916 509134
rect 163152 508898 168847 509134
rect 169083 508898 190916 509134
rect 191152 508898 196847 509134
rect 197083 508898 218916 509134
rect 219152 508898 224847 509134
rect 225083 508898 246916 509134
rect 247152 508898 252847 509134
rect 253083 508898 274916 509134
rect 275152 508898 280847 509134
rect 281083 508898 302916 509134
rect 303152 508898 308847 509134
rect 309083 508898 330916 509134
rect 331152 508898 336847 509134
rect 337083 508898 358916 509134
rect 359152 508898 364847 509134
rect 365083 508898 386916 509134
rect 387152 508898 392847 509134
rect 393083 508898 414916 509134
rect 415152 508898 420847 509134
rect 421083 508898 442916 509134
rect 443152 508898 448847 509134
rect 449083 508898 470916 509134
rect 471152 508898 476847 509134
rect 477083 508898 498916 509134
rect 499152 508898 504847 509134
rect 505083 508898 526916 509134
rect 527152 508898 532847 509134
rect 533083 508898 554916 509134
rect 555152 508898 560847 509134
rect 561083 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 592650 509134
rect -8726 508866 592650 508898
rect -8726 485829 592650 485861
rect -8726 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 19952 485829
rect 20188 485593 25882 485829
rect 26118 485593 31813 485829
rect 32049 485593 47952 485829
rect 48188 485593 53882 485829
rect 54118 485593 59813 485829
rect 60049 485593 75952 485829
rect 76188 485593 81882 485829
rect 82118 485593 87813 485829
rect 88049 485593 103952 485829
rect 104188 485593 109882 485829
rect 110118 485593 115813 485829
rect 116049 485593 131952 485829
rect 132188 485593 137882 485829
rect 138118 485593 143813 485829
rect 144049 485593 159952 485829
rect 160188 485593 165882 485829
rect 166118 485593 171813 485829
rect 172049 485593 187952 485829
rect 188188 485593 193882 485829
rect 194118 485593 199813 485829
rect 200049 485593 215952 485829
rect 216188 485593 221882 485829
rect 222118 485593 227813 485829
rect 228049 485593 243952 485829
rect 244188 485593 249882 485829
rect 250118 485593 255813 485829
rect 256049 485593 271952 485829
rect 272188 485593 277882 485829
rect 278118 485593 283813 485829
rect 284049 485593 299952 485829
rect 300188 485593 305882 485829
rect 306118 485593 311813 485829
rect 312049 485593 327952 485829
rect 328188 485593 333882 485829
rect 334118 485593 339813 485829
rect 340049 485593 355952 485829
rect 356188 485593 361882 485829
rect 362118 485593 367813 485829
rect 368049 485593 383952 485829
rect 384188 485593 389882 485829
rect 390118 485593 395813 485829
rect 396049 485593 411952 485829
rect 412188 485593 417882 485829
rect 418118 485593 423813 485829
rect 424049 485593 439952 485829
rect 440188 485593 445882 485829
rect 446118 485593 451813 485829
rect 452049 485593 467952 485829
rect 468188 485593 473882 485829
rect 474118 485593 479813 485829
rect 480049 485593 495952 485829
rect 496188 485593 501882 485829
rect 502118 485593 507813 485829
rect 508049 485593 523952 485829
rect 524188 485593 529882 485829
rect 530118 485593 535813 485829
rect 536049 485593 551952 485829
rect 552188 485593 557882 485829
rect 558118 485593 563813 485829
rect 564049 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 592650 485829
rect -8726 485509 592650 485593
rect -8726 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 19952 485509
rect 20188 485273 25882 485509
rect 26118 485273 31813 485509
rect 32049 485273 47952 485509
rect 48188 485273 53882 485509
rect 54118 485273 59813 485509
rect 60049 485273 75952 485509
rect 76188 485273 81882 485509
rect 82118 485273 87813 485509
rect 88049 485273 103952 485509
rect 104188 485273 109882 485509
rect 110118 485273 115813 485509
rect 116049 485273 131952 485509
rect 132188 485273 137882 485509
rect 138118 485273 143813 485509
rect 144049 485273 159952 485509
rect 160188 485273 165882 485509
rect 166118 485273 171813 485509
rect 172049 485273 187952 485509
rect 188188 485273 193882 485509
rect 194118 485273 199813 485509
rect 200049 485273 215952 485509
rect 216188 485273 221882 485509
rect 222118 485273 227813 485509
rect 228049 485273 243952 485509
rect 244188 485273 249882 485509
rect 250118 485273 255813 485509
rect 256049 485273 271952 485509
rect 272188 485273 277882 485509
rect 278118 485273 283813 485509
rect 284049 485273 299952 485509
rect 300188 485273 305882 485509
rect 306118 485273 311813 485509
rect 312049 485273 327952 485509
rect 328188 485273 333882 485509
rect 334118 485273 339813 485509
rect 340049 485273 355952 485509
rect 356188 485273 361882 485509
rect 362118 485273 367813 485509
rect 368049 485273 383952 485509
rect 384188 485273 389882 485509
rect 390118 485273 395813 485509
rect 396049 485273 411952 485509
rect 412188 485273 417882 485509
rect 418118 485273 423813 485509
rect 424049 485273 439952 485509
rect 440188 485273 445882 485509
rect 446118 485273 451813 485509
rect 452049 485273 467952 485509
rect 468188 485273 473882 485509
rect 474118 485273 479813 485509
rect 480049 485273 495952 485509
rect 496188 485273 501882 485509
rect 502118 485273 507813 485509
rect 508049 485273 523952 485509
rect 524188 485273 529882 485509
rect 530118 485273 535813 485509
rect 536049 485273 551952 485509
rect 552188 485273 557882 485509
rect 558118 485273 563813 485509
rect 564049 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 592650 485509
rect -8726 485241 592650 485273
rect -8726 482454 592650 482486
rect -8726 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 22916 482454
rect 23152 482218 28847 482454
rect 29083 482218 50916 482454
rect 51152 482218 56847 482454
rect 57083 482218 78916 482454
rect 79152 482218 84847 482454
rect 85083 482218 106916 482454
rect 107152 482218 112847 482454
rect 113083 482218 134916 482454
rect 135152 482218 140847 482454
rect 141083 482218 162916 482454
rect 163152 482218 168847 482454
rect 169083 482218 190916 482454
rect 191152 482218 196847 482454
rect 197083 482218 218916 482454
rect 219152 482218 224847 482454
rect 225083 482218 246916 482454
rect 247152 482218 252847 482454
rect 253083 482218 274916 482454
rect 275152 482218 280847 482454
rect 281083 482218 302916 482454
rect 303152 482218 308847 482454
rect 309083 482218 330916 482454
rect 331152 482218 336847 482454
rect 337083 482218 358916 482454
rect 359152 482218 364847 482454
rect 365083 482218 386916 482454
rect 387152 482218 392847 482454
rect 393083 482218 414916 482454
rect 415152 482218 420847 482454
rect 421083 482218 442916 482454
rect 443152 482218 448847 482454
rect 449083 482218 470916 482454
rect 471152 482218 476847 482454
rect 477083 482218 498916 482454
rect 499152 482218 504847 482454
rect 505083 482218 526916 482454
rect 527152 482218 532847 482454
rect 533083 482218 554916 482454
rect 555152 482218 560847 482454
rect 561083 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 592650 482454
rect -8726 482134 592650 482218
rect -8726 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 22916 482134
rect 23152 481898 28847 482134
rect 29083 481898 50916 482134
rect 51152 481898 56847 482134
rect 57083 481898 78916 482134
rect 79152 481898 84847 482134
rect 85083 481898 106916 482134
rect 107152 481898 112847 482134
rect 113083 481898 134916 482134
rect 135152 481898 140847 482134
rect 141083 481898 162916 482134
rect 163152 481898 168847 482134
rect 169083 481898 190916 482134
rect 191152 481898 196847 482134
rect 197083 481898 218916 482134
rect 219152 481898 224847 482134
rect 225083 481898 246916 482134
rect 247152 481898 252847 482134
rect 253083 481898 274916 482134
rect 275152 481898 280847 482134
rect 281083 481898 302916 482134
rect 303152 481898 308847 482134
rect 309083 481898 330916 482134
rect 331152 481898 336847 482134
rect 337083 481898 358916 482134
rect 359152 481898 364847 482134
rect 365083 481898 386916 482134
rect 387152 481898 392847 482134
rect 393083 481898 414916 482134
rect 415152 481898 420847 482134
rect 421083 481898 442916 482134
rect 443152 481898 448847 482134
rect 449083 481898 470916 482134
rect 471152 481898 476847 482134
rect 477083 481898 498916 482134
rect 499152 481898 504847 482134
rect 505083 481898 526916 482134
rect 527152 481898 532847 482134
rect 533083 481898 554916 482134
rect 555152 481898 560847 482134
rect 561083 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 592650 482134
rect -8726 481866 592650 481898
rect -8726 458829 592650 458861
rect -8726 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 19952 458829
rect 20188 458593 25882 458829
rect 26118 458593 31813 458829
rect 32049 458593 47952 458829
rect 48188 458593 53882 458829
rect 54118 458593 59813 458829
rect 60049 458593 75952 458829
rect 76188 458593 81882 458829
rect 82118 458593 87813 458829
rect 88049 458593 103952 458829
rect 104188 458593 109882 458829
rect 110118 458593 115813 458829
rect 116049 458593 131952 458829
rect 132188 458593 137882 458829
rect 138118 458593 143813 458829
rect 144049 458593 159952 458829
rect 160188 458593 165882 458829
rect 166118 458593 171813 458829
rect 172049 458593 187952 458829
rect 188188 458593 193882 458829
rect 194118 458593 199813 458829
rect 200049 458593 215952 458829
rect 216188 458593 221882 458829
rect 222118 458593 227813 458829
rect 228049 458593 243952 458829
rect 244188 458593 249882 458829
rect 250118 458593 255813 458829
rect 256049 458593 271952 458829
rect 272188 458593 277882 458829
rect 278118 458593 283813 458829
rect 284049 458593 299952 458829
rect 300188 458593 305882 458829
rect 306118 458593 311813 458829
rect 312049 458593 327952 458829
rect 328188 458593 333882 458829
rect 334118 458593 339813 458829
rect 340049 458593 355952 458829
rect 356188 458593 361882 458829
rect 362118 458593 367813 458829
rect 368049 458593 383952 458829
rect 384188 458593 389882 458829
rect 390118 458593 395813 458829
rect 396049 458593 411952 458829
rect 412188 458593 417882 458829
rect 418118 458593 423813 458829
rect 424049 458593 439952 458829
rect 440188 458593 445882 458829
rect 446118 458593 451813 458829
rect 452049 458593 467952 458829
rect 468188 458593 473882 458829
rect 474118 458593 479813 458829
rect 480049 458593 495952 458829
rect 496188 458593 501882 458829
rect 502118 458593 507813 458829
rect 508049 458593 523952 458829
rect 524188 458593 529882 458829
rect 530118 458593 535813 458829
rect 536049 458593 551952 458829
rect 552188 458593 557882 458829
rect 558118 458593 563813 458829
rect 564049 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 592650 458829
rect -8726 458509 592650 458593
rect -8726 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 19952 458509
rect 20188 458273 25882 458509
rect 26118 458273 31813 458509
rect 32049 458273 47952 458509
rect 48188 458273 53882 458509
rect 54118 458273 59813 458509
rect 60049 458273 75952 458509
rect 76188 458273 81882 458509
rect 82118 458273 87813 458509
rect 88049 458273 103952 458509
rect 104188 458273 109882 458509
rect 110118 458273 115813 458509
rect 116049 458273 131952 458509
rect 132188 458273 137882 458509
rect 138118 458273 143813 458509
rect 144049 458273 159952 458509
rect 160188 458273 165882 458509
rect 166118 458273 171813 458509
rect 172049 458273 187952 458509
rect 188188 458273 193882 458509
rect 194118 458273 199813 458509
rect 200049 458273 215952 458509
rect 216188 458273 221882 458509
rect 222118 458273 227813 458509
rect 228049 458273 243952 458509
rect 244188 458273 249882 458509
rect 250118 458273 255813 458509
rect 256049 458273 271952 458509
rect 272188 458273 277882 458509
rect 278118 458273 283813 458509
rect 284049 458273 299952 458509
rect 300188 458273 305882 458509
rect 306118 458273 311813 458509
rect 312049 458273 327952 458509
rect 328188 458273 333882 458509
rect 334118 458273 339813 458509
rect 340049 458273 355952 458509
rect 356188 458273 361882 458509
rect 362118 458273 367813 458509
rect 368049 458273 383952 458509
rect 384188 458273 389882 458509
rect 390118 458273 395813 458509
rect 396049 458273 411952 458509
rect 412188 458273 417882 458509
rect 418118 458273 423813 458509
rect 424049 458273 439952 458509
rect 440188 458273 445882 458509
rect 446118 458273 451813 458509
rect 452049 458273 467952 458509
rect 468188 458273 473882 458509
rect 474118 458273 479813 458509
rect 480049 458273 495952 458509
rect 496188 458273 501882 458509
rect 502118 458273 507813 458509
rect 508049 458273 523952 458509
rect 524188 458273 529882 458509
rect 530118 458273 535813 458509
rect 536049 458273 551952 458509
rect 552188 458273 557882 458509
rect 558118 458273 563813 458509
rect 564049 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 592650 458509
rect -8726 458241 592650 458273
rect -8726 455454 592650 455486
rect -8726 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 22916 455454
rect 23152 455218 28847 455454
rect 29083 455218 50916 455454
rect 51152 455218 56847 455454
rect 57083 455218 78916 455454
rect 79152 455218 84847 455454
rect 85083 455218 106916 455454
rect 107152 455218 112847 455454
rect 113083 455218 134916 455454
rect 135152 455218 140847 455454
rect 141083 455218 162916 455454
rect 163152 455218 168847 455454
rect 169083 455218 190916 455454
rect 191152 455218 196847 455454
rect 197083 455218 218916 455454
rect 219152 455218 224847 455454
rect 225083 455218 246916 455454
rect 247152 455218 252847 455454
rect 253083 455218 274916 455454
rect 275152 455218 280847 455454
rect 281083 455218 302916 455454
rect 303152 455218 308847 455454
rect 309083 455218 330916 455454
rect 331152 455218 336847 455454
rect 337083 455218 358916 455454
rect 359152 455218 364847 455454
rect 365083 455218 386916 455454
rect 387152 455218 392847 455454
rect 393083 455218 414916 455454
rect 415152 455218 420847 455454
rect 421083 455218 442916 455454
rect 443152 455218 448847 455454
rect 449083 455218 470916 455454
rect 471152 455218 476847 455454
rect 477083 455218 498916 455454
rect 499152 455218 504847 455454
rect 505083 455218 526916 455454
rect 527152 455218 532847 455454
rect 533083 455218 554916 455454
rect 555152 455218 560847 455454
rect 561083 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 592650 455454
rect -8726 455134 592650 455218
rect -8726 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 22916 455134
rect 23152 454898 28847 455134
rect 29083 454898 50916 455134
rect 51152 454898 56847 455134
rect 57083 454898 78916 455134
rect 79152 454898 84847 455134
rect 85083 454898 106916 455134
rect 107152 454898 112847 455134
rect 113083 454898 134916 455134
rect 135152 454898 140847 455134
rect 141083 454898 162916 455134
rect 163152 454898 168847 455134
rect 169083 454898 190916 455134
rect 191152 454898 196847 455134
rect 197083 454898 218916 455134
rect 219152 454898 224847 455134
rect 225083 454898 246916 455134
rect 247152 454898 252847 455134
rect 253083 454898 274916 455134
rect 275152 454898 280847 455134
rect 281083 454898 302916 455134
rect 303152 454898 308847 455134
rect 309083 454898 330916 455134
rect 331152 454898 336847 455134
rect 337083 454898 358916 455134
rect 359152 454898 364847 455134
rect 365083 454898 386916 455134
rect 387152 454898 392847 455134
rect 393083 454898 414916 455134
rect 415152 454898 420847 455134
rect 421083 454898 442916 455134
rect 443152 454898 448847 455134
rect 449083 454898 470916 455134
rect 471152 454898 476847 455134
rect 477083 454898 498916 455134
rect 499152 454898 504847 455134
rect 505083 454898 526916 455134
rect 527152 454898 532847 455134
rect 533083 454898 554916 455134
rect 555152 454898 560847 455134
rect 561083 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 592650 455134
rect -8726 454866 592650 454898
rect -8726 431829 592650 431861
rect -8726 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 19952 431829
rect 20188 431593 25882 431829
rect 26118 431593 31813 431829
rect 32049 431593 47952 431829
rect 48188 431593 53882 431829
rect 54118 431593 59813 431829
rect 60049 431593 75952 431829
rect 76188 431593 81882 431829
rect 82118 431593 87813 431829
rect 88049 431593 103952 431829
rect 104188 431593 109882 431829
rect 110118 431593 115813 431829
rect 116049 431593 131952 431829
rect 132188 431593 137882 431829
rect 138118 431593 143813 431829
rect 144049 431593 159952 431829
rect 160188 431593 165882 431829
rect 166118 431593 171813 431829
rect 172049 431593 187952 431829
rect 188188 431593 193882 431829
rect 194118 431593 199813 431829
rect 200049 431593 215952 431829
rect 216188 431593 221882 431829
rect 222118 431593 227813 431829
rect 228049 431593 243952 431829
rect 244188 431593 249882 431829
rect 250118 431593 255813 431829
rect 256049 431593 271952 431829
rect 272188 431593 277882 431829
rect 278118 431593 283813 431829
rect 284049 431593 299952 431829
rect 300188 431593 305882 431829
rect 306118 431593 311813 431829
rect 312049 431593 327952 431829
rect 328188 431593 333882 431829
rect 334118 431593 339813 431829
rect 340049 431593 355952 431829
rect 356188 431593 361882 431829
rect 362118 431593 367813 431829
rect 368049 431593 383952 431829
rect 384188 431593 389882 431829
rect 390118 431593 395813 431829
rect 396049 431593 411952 431829
rect 412188 431593 417882 431829
rect 418118 431593 423813 431829
rect 424049 431593 439952 431829
rect 440188 431593 445882 431829
rect 446118 431593 451813 431829
rect 452049 431593 467952 431829
rect 468188 431593 473882 431829
rect 474118 431593 479813 431829
rect 480049 431593 495952 431829
rect 496188 431593 501882 431829
rect 502118 431593 507813 431829
rect 508049 431593 523952 431829
rect 524188 431593 529882 431829
rect 530118 431593 535813 431829
rect 536049 431593 551952 431829
rect 552188 431593 557882 431829
rect 558118 431593 563813 431829
rect 564049 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 592650 431829
rect -8726 431509 592650 431593
rect -8726 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 19952 431509
rect 20188 431273 25882 431509
rect 26118 431273 31813 431509
rect 32049 431273 47952 431509
rect 48188 431273 53882 431509
rect 54118 431273 59813 431509
rect 60049 431273 75952 431509
rect 76188 431273 81882 431509
rect 82118 431273 87813 431509
rect 88049 431273 103952 431509
rect 104188 431273 109882 431509
rect 110118 431273 115813 431509
rect 116049 431273 131952 431509
rect 132188 431273 137882 431509
rect 138118 431273 143813 431509
rect 144049 431273 159952 431509
rect 160188 431273 165882 431509
rect 166118 431273 171813 431509
rect 172049 431273 187952 431509
rect 188188 431273 193882 431509
rect 194118 431273 199813 431509
rect 200049 431273 215952 431509
rect 216188 431273 221882 431509
rect 222118 431273 227813 431509
rect 228049 431273 243952 431509
rect 244188 431273 249882 431509
rect 250118 431273 255813 431509
rect 256049 431273 271952 431509
rect 272188 431273 277882 431509
rect 278118 431273 283813 431509
rect 284049 431273 299952 431509
rect 300188 431273 305882 431509
rect 306118 431273 311813 431509
rect 312049 431273 327952 431509
rect 328188 431273 333882 431509
rect 334118 431273 339813 431509
rect 340049 431273 355952 431509
rect 356188 431273 361882 431509
rect 362118 431273 367813 431509
rect 368049 431273 383952 431509
rect 384188 431273 389882 431509
rect 390118 431273 395813 431509
rect 396049 431273 411952 431509
rect 412188 431273 417882 431509
rect 418118 431273 423813 431509
rect 424049 431273 439952 431509
rect 440188 431273 445882 431509
rect 446118 431273 451813 431509
rect 452049 431273 467952 431509
rect 468188 431273 473882 431509
rect 474118 431273 479813 431509
rect 480049 431273 495952 431509
rect 496188 431273 501882 431509
rect 502118 431273 507813 431509
rect 508049 431273 523952 431509
rect 524188 431273 529882 431509
rect 530118 431273 535813 431509
rect 536049 431273 551952 431509
rect 552188 431273 557882 431509
rect 558118 431273 563813 431509
rect 564049 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 592650 431509
rect -8726 431241 592650 431273
rect -8726 428454 592650 428486
rect -8726 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 22916 428454
rect 23152 428218 28847 428454
rect 29083 428218 50916 428454
rect 51152 428218 56847 428454
rect 57083 428218 78916 428454
rect 79152 428218 84847 428454
rect 85083 428218 106916 428454
rect 107152 428218 112847 428454
rect 113083 428218 134916 428454
rect 135152 428218 140847 428454
rect 141083 428218 162916 428454
rect 163152 428218 168847 428454
rect 169083 428218 190916 428454
rect 191152 428218 196847 428454
rect 197083 428218 218916 428454
rect 219152 428218 224847 428454
rect 225083 428218 246916 428454
rect 247152 428218 252847 428454
rect 253083 428218 274916 428454
rect 275152 428218 280847 428454
rect 281083 428218 302916 428454
rect 303152 428218 308847 428454
rect 309083 428218 330916 428454
rect 331152 428218 336847 428454
rect 337083 428218 358916 428454
rect 359152 428218 364847 428454
rect 365083 428218 386916 428454
rect 387152 428218 392847 428454
rect 393083 428218 414916 428454
rect 415152 428218 420847 428454
rect 421083 428218 442916 428454
rect 443152 428218 448847 428454
rect 449083 428218 470916 428454
rect 471152 428218 476847 428454
rect 477083 428218 498916 428454
rect 499152 428218 504847 428454
rect 505083 428218 526916 428454
rect 527152 428218 532847 428454
rect 533083 428218 554916 428454
rect 555152 428218 560847 428454
rect 561083 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 592650 428454
rect -8726 428134 592650 428218
rect -8726 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 22916 428134
rect 23152 427898 28847 428134
rect 29083 427898 50916 428134
rect 51152 427898 56847 428134
rect 57083 427898 78916 428134
rect 79152 427898 84847 428134
rect 85083 427898 106916 428134
rect 107152 427898 112847 428134
rect 113083 427898 134916 428134
rect 135152 427898 140847 428134
rect 141083 427898 162916 428134
rect 163152 427898 168847 428134
rect 169083 427898 190916 428134
rect 191152 427898 196847 428134
rect 197083 427898 218916 428134
rect 219152 427898 224847 428134
rect 225083 427898 246916 428134
rect 247152 427898 252847 428134
rect 253083 427898 274916 428134
rect 275152 427898 280847 428134
rect 281083 427898 302916 428134
rect 303152 427898 308847 428134
rect 309083 427898 330916 428134
rect 331152 427898 336847 428134
rect 337083 427898 358916 428134
rect 359152 427898 364847 428134
rect 365083 427898 386916 428134
rect 387152 427898 392847 428134
rect 393083 427898 414916 428134
rect 415152 427898 420847 428134
rect 421083 427898 442916 428134
rect 443152 427898 448847 428134
rect 449083 427898 470916 428134
rect 471152 427898 476847 428134
rect 477083 427898 498916 428134
rect 499152 427898 504847 428134
rect 505083 427898 526916 428134
rect 527152 427898 532847 428134
rect 533083 427898 554916 428134
rect 555152 427898 560847 428134
rect 561083 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 592650 428134
rect -8726 427866 592650 427898
rect -8726 404829 592650 404861
rect -8726 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 19952 404829
rect 20188 404593 25882 404829
rect 26118 404593 31813 404829
rect 32049 404593 47952 404829
rect 48188 404593 53882 404829
rect 54118 404593 59813 404829
rect 60049 404593 75952 404829
rect 76188 404593 81882 404829
rect 82118 404593 87813 404829
rect 88049 404593 103952 404829
rect 104188 404593 109882 404829
rect 110118 404593 115813 404829
rect 116049 404593 131952 404829
rect 132188 404593 137882 404829
rect 138118 404593 143813 404829
rect 144049 404593 159952 404829
rect 160188 404593 165882 404829
rect 166118 404593 171813 404829
rect 172049 404593 187952 404829
rect 188188 404593 193882 404829
rect 194118 404593 199813 404829
rect 200049 404593 215952 404829
rect 216188 404593 221882 404829
rect 222118 404593 227813 404829
rect 228049 404593 243952 404829
rect 244188 404593 249882 404829
rect 250118 404593 255813 404829
rect 256049 404593 271952 404829
rect 272188 404593 277882 404829
rect 278118 404593 283813 404829
rect 284049 404593 299952 404829
rect 300188 404593 305882 404829
rect 306118 404593 311813 404829
rect 312049 404593 327952 404829
rect 328188 404593 333882 404829
rect 334118 404593 339813 404829
rect 340049 404593 355952 404829
rect 356188 404593 361882 404829
rect 362118 404593 367813 404829
rect 368049 404593 383952 404829
rect 384188 404593 389882 404829
rect 390118 404593 395813 404829
rect 396049 404593 411952 404829
rect 412188 404593 417882 404829
rect 418118 404593 423813 404829
rect 424049 404593 439952 404829
rect 440188 404593 445882 404829
rect 446118 404593 451813 404829
rect 452049 404593 467952 404829
rect 468188 404593 473882 404829
rect 474118 404593 479813 404829
rect 480049 404593 495952 404829
rect 496188 404593 501882 404829
rect 502118 404593 507813 404829
rect 508049 404593 523952 404829
rect 524188 404593 529882 404829
rect 530118 404593 535813 404829
rect 536049 404593 551952 404829
rect 552188 404593 557882 404829
rect 558118 404593 563813 404829
rect 564049 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 592650 404829
rect -8726 404509 592650 404593
rect -8726 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 19952 404509
rect 20188 404273 25882 404509
rect 26118 404273 31813 404509
rect 32049 404273 47952 404509
rect 48188 404273 53882 404509
rect 54118 404273 59813 404509
rect 60049 404273 75952 404509
rect 76188 404273 81882 404509
rect 82118 404273 87813 404509
rect 88049 404273 103952 404509
rect 104188 404273 109882 404509
rect 110118 404273 115813 404509
rect 116049 404273 131952 404509
rect 132188 404273 137882 404509
rect 138118 404273 143813 404509
rect 144049 404273 159952 404509
rect 160188 404273 165882 404509
rect 166118 404273 171813 404509
rect 172049 404273 187952 404509
rect 188188 404273 193882 404509
rect 194118 404273 199813 404509
rect 200049 404273 215952 404509
rect 216188 404273 221882 404509
rect 222118 404273 227813 404509
rect 228049 404273 243952 404509
rect 244188 404273 249882 404509
rect 250118 404273 255813 404509
rect 256049 404273 271952 404509
rect 272188 404273 277882 404509
rect 278118 404273 283813 404509
rect 284049 404273 299952 404509
rect 300188 404273 305882 404509
rect 306118 404273 311813 404509
rect 312049 404273 327952 404509
rect 328188 404273 333882 404509
rect 334118 404273 339813 404509
rect 340049 404273 355952 404509
rect 356188 404273 361882 404509
rect 362118 404273 367813 404509
rect 368049 404273 383952 404509
rect 384188 404273 389882 404509
rect 390118 404273 395813 404509
rect 396049 404273 411952 404509
rect 412188 404273 417882 404509
rect 418118 404273 423813 404509
rect 424049 404273 439952 404509
rect 440188 404273 445882 404509
rect 446118 404273 451813 404509
rect 452049 404273 467952 404509
rect 468188 404273 473882 404509
rect 474118 404273 479813 404509
rect 480049 404273 495952 404509
rect 496188 404273 501882 404509
rect 502118 404273 507813 404509
rect 508049 404273 523952 404509
rect 524188 404273 529882 404509
rect 530118 404273 535813 404509
rect 536049 404273 551952 404509
rect 552188 404273 557882 404509
rect 558118 404273 563813 404509
rect 564049 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 592650 404509
rect -8726 404241 592650 404273
rect -8726 401454 592650 401486
rect -8726 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 22916 401454
rect 23152 401218 28847 401454
rect 29083 401218 50916 401454
rect 51152 401218 56847 401454
rect 57083 401218 78916 401454
rect 79152 401218 84847 401454
rect 85083 401218 106916 401454
rect 107152 401218 112847 401454
rect 113083 401218 134916 401454
rect 135152 401218 140847 401454
rect 141083 401218 162916 401454
rect 163152 401218 168847 401454
rect 169083 401218 190916 401454
rect 191152 401218 196847 401454
rect 197083 401218 218916 401454
rect 219152 401218 224847 401454
rect 225083 401218 246916 401454
rect 247152 401218 252847 401454
rect 253083 401218 274916 401454
rect 275152 401218 280847 401454
rect 281083 401218 302916 401454
rect 303152 401218 308847 401454
rect 309083 401218 330916 401454
rect 331152 401218 336847 401454
rect 337083 401218 358916 401454
rect 359152 401218 364847 401454
rect 365083 401218 386916 401454
rect 387152 401218 392847 401454
rect 393083 401218 414916 401454
rect 415152 401218 420847 401454
rect 421083 401218 442916 401454
rect 443152 401218 448847 401454
rect 449083 401218 470916 401454
rect 471152 401218 476847 401454
rect 477083 401218 498916 401454
rect 499152 401218 504847 401454
rect 505083 401218 526916 401454
rect 527152 401218 532847 401454
rect 533083 401218 554916 401454
rect 555152 401218 560847 401454
rect 561083 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 592650 401454
rect -8726 401134 592650 401218
rect -8726 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 22916 401134
rect 23152 400898 28847 401134
rect 29083 400898 50916 401134
rect 51152 400898 56847 401134
rect 57083 400898 78916 401134
rect 79152 400898 84847 401134
rect 85083 400898 106916 401134
rect 107152 400898 112847 401134
rect 113083 400898 134916 401134
rect 135152 400898 140847 401134
rect 141083 400898 162916 401134
rect 163152 400898 168847 401134
rect 169083 400898 190916 401134
rect 191152 400898 196847 401134
rect 197083 400898 218916 401134
rect 219152 400898 224847 401134
rect 225083 400898 246916 401134
rect 247152 400898 252847 401134
rect 253083 400898 274916 401134
rect 275152 400898 280847 401134
rect 281083 400898 302916 401134
rect 303152 400898 308847 401134
rect 309083 400898 330916 401134
rect 331152 400898 336847 401134
rect 337083 400898 358916 401134
rect 359152 400898 364847 401134
rect 365083 400898 386916 401134
rect 387152 400898 392847 401134
rect 393083 400898 414916 401134
rect 415152 400898 420847 401134
rect 421083 400898 442916 401134
rect 443152 400898 448847 401134
rect 449083 400898 470916 401134
rect 471152 400898 476847 401134
rect 477083 400898 498916 401134
rect 499152 400898 504847 401134
rect 505083 400898 526916 401134
rect 527152 400898 532847 401134
rect 533083 400898 554916 401134
rect 555152 400898 560847 401134
rect 561083 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 592650 401134
rect -8726 400866 592650 400898
rect -8726 377829 592650 377861
rect -8726 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 19952 377829
rect 20188 377593 25882 377829
rect 26118 377593 31813 377829
rect 32049 377593 47952 377829
rect 48188 377593 53882 377829
rect 54118 377593 59813 377829
rect 60049 377593 75952 377829
rect 76188 377593 81882 377829
rect 82118 377593 87813 377829
rect 88049 377593 103952 377829
rect 104188 377593 109882 377829
rect 110118 377593 115813 377829
rect 116049 377593 131952 377829
rect 132188 377593 137882 377829
rect 138118 377593 143813 377829
rect 144049 377593 159952 377829
rect 160188 377593 165882 377829
rect 166118 377593 171813 377829
rect 172049 377593 187952 377829
rect 188188 377593 193882 377829
rect 194118 377593 199813 377829
rect 200049 377593 215952 377829
rect 216188 377593 221882 377829
rect 222118 377593 227813 377829
rect 228049 377593 243952 377829
rect 244188 377593 249882 377829
rect 250118 377593 255813 377829
rect 256049 377593 271952 377829
rect 272188 377593 277882 377829
rect 278118 377593 283813 377829
rect 284049 377593 299952 377829
rect 300188 377593 305882 377829
rect 306118 377593 311813 377829
rect 312049 377593 327952 377829
rect 328188 377593 333882 377829
rect 334118 377593 339813 377829
rect 340049 377593 355952 377829
rect 356188 377593 361882 377829
rect 362118 377593 367813 377829
rect 368049 377593 383952 377829
rect 384188 377593 389882 377829
rect 390118 377593 395813 377829
rect 396049 377593 411952 377829
rect 412188 377593 417882 377829
rect 418118 377593 423813 377829
rect 424049 377593 439952 377829
rect 440188 377593 445882 377829
rect 446118 377593 451813 377829
rect 452049 377593 467952 377829
rect 468188 377593 473882 377829
rect 474118 377593 479813 377829
rect 480049 377593 495952 377829
rect 496188 377593 501882 377829
rect 502118 377593 507813 377829
rect 508049 377593 523952 377829
rect 524188 377593 529882 377829
rect 530118 377593 535813 377829
rect 536049 377593 551952 377829
rect 552188 377593 557882 377829
rect 558118 377593 563813 377829
rect 564049 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 592650 377829
rect -8726 377509 592650 377593
rect -8726 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 19952 377509
rect 20188 377273 25882 377509
rect 26118 377273 31813 377509
rect 32049 377273 47952 377509
rect 48188 377273 53882 377509
rect 54118 377273 59813 377509
rect 60049 377273 75952 377509
rect 76188 377273 81882 377509
rect 82118 377273 87813 377509
rect 88049 377273 103952 377509
rect 104188 377273 109882 377509
rect 110118 377273 115813 377509
rect 116049 377273 131952 377509
rect 132188 377273 137882 377509
rect 138118 377273 143813 377509
rect 144049 377273 159952 377509
rect 160188 377273 165882 377509
rect 166118 377273 171813 377509
rect 172049 377273 187952 377509
rect 188188 377273 193882 377509
rect 194118 377273 199813 377509
rect 200049 377273 215952 377509
rect 216188 377273 221882 377509
rect 222118 377273 227813 377509
rect 228049 377273 243952 377509
rect 244188 377273 249882 377509
rect 250118 377273 255813 377509
rect 256049 377273 271952 377509
rect 272188 377273 277882 377509
rect 278118 377273 283813 377509
rect 284049 377273 299952 377509
rect 300188 377273 305882 377509
rect 306118 377273 311813 377509
rect 312049 377273 327952 377509
rect 328188 377273 333882 377509
rect 334118 377273 339813 377509
rect 340049 377273 355952 377509
rect 356188 377273 361882 377509
rect 362118 377273 367813 377509
rect 368049 377273 383952 377509
rect 384188 377273 389882 377509
rect 390118 377273 395813 377509
rect 396049 377273 411952 377509
rect 412188 377273 417882 377509
rect 418118 377273 423813 377509
rect 424049 377273 439952 377509
rect 440188 377273 445882 377509
rect 446118 377273 451813 377509
rect 452049 377273 467952 377509
rect 468188 377273 473882 377509
rect 474118 377273 479813 377509
rect 480049 377273 495952 377509
rect 496188 377273 501882 377509
rect 502118 377273 507813 377509
rect 508049 377273 523952 377509
rect 524188 377273 529882 377509
rect 530118 377273 535813 377509
rect 536049 377273 551952 377509
rect 552188 377273 557882 377509
rect 558118 377273 563813 377509
rect 564049 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 592650 377509
rect -8726 377241 592650 377273
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 22916 374454
rect 23152 374218 28847 374454
rect 29083 374218 50916 374454
rect 51152 374218 56847 374454
rect 57083 374218 78916 374454
rect 79152 374218 84847 374454
rect 85083 374218 106916 374454
rect 107152 374218 112847 374454
rect 113083 374218 134916 374454
rect 135152 374218 140847 374454
rect 141083 374218 162916 374454
rect 163152 374218 168847 374454
rect 169083 374218 190916 374454
rect 191152 374218 196847 374454
rect 197083 374218 218916 374454
rect 219152 374218 224847 374454
rect 225083 374218 246916 374454
rect 247152 374218 252847 374454
rect 253083 374218 274916 374454
rect 275152 374218 280847 374454
rect 281083 374218 302916 374454
rect 303152 374218 308847 374454
rect 309083 374218 330916 374454
rect 331152 374218 336847 374454
rect 337083 374218 358916 374454
rect 359152 374218 364847 374454
rect 365083 374218 386916 374454
rect 387152 374218 392847 374454
rect 393083 374218 414916 374454
rect 415152 374218 420847 374454
rect 421083 374218 442916 374454
rect 443152 374218 448847 374454
rect 449083 374218 470916 374454
rect 471152 374218 476847 374454
rect 477083 374218 498916 374454
rect 499152 374218 504847 374454
rect 505083 374218 526916 374454
rect 527152 374218 532847 374454
rect 533083 374218 554916 374454
rect 555152 374218 560847 374454
rect 561083 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 22916 374134
rect 23152 373898 28847 374134
rect 29083 373898 50916 374134
rect 51152 373898 56847 374134
rect 57083 373898 78916 374134
rect 79152 373898 84847 374134
rect 85083 373898 106916 374134
rect 107152 373898 112847 374134
rect 113083 373898 134916 374134
rect 135152 373898 140847 374134
rect 141083 373898 162916 374134
rect 163152 373898 168847 374134
rect 169083 373898 190916 374134
rect 191152 373898 196847 374134
rect 197083 373898 218916 374134
rect 219152 373898 224847 374134
rect 225083 373898 246916 374134
rect 247152 373898 252847 374134
rect 253083 373898 274916 374134
rect 275152 373898 280847 374134
rect 281083 373898 302916 374134
rect 303152 373898 308847 374134
rect 309083 373898 330916 374134
rect 331152 373898 336847 374134
rect 337083 373898 358916 374134
rect 359152 373898 364847 374134
rect 365083 373898 386916 374134
rect 387152 373898 392847 374134
rect 393083 373898 414916 374134
rect 415152 373898 420847 374134
rect 421083 373898 442916 374134
rect 443152 373898 448847 374134
rect 449083 373898 470916 374134
rect 471152 373898 476847 374134
rect 477083 373898 498916 374134
rect 499152 373898 504847 374134
rect 505083 373898 526916 374134
rect 527152 373898 532847 374134
rect 533083 373898 554916 374134
rect 555152 373898 560847 374134
rect 561083 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 350829 592650 350861
rect -8726 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 19952 350829
rect 20188 350593 25882 350829
rect 26118 350593 31813 350829
rect 32049 350593 47952 350829
rect 48188 350593 53882 350829
rect 54118 350593 59813 350829
rect 60049 350593 75952 350829
rect 76188 350593 81882 350829
rect 82118 350593 87813 350829
rect 88049 350593 103952 350829
rect 104188 350593 109882 350829
rect 110118 350593 115813 350829
rect 116049 350593 131952 350829
rect 132188 350593 137882 350829
rect 138118 350593 143813 350829
rect 144049 350593 159952 350829
rect 160188 350593 165882 350829
rect 166118 350593 171813 350829
rect 172049 350593 187952 350829
rect 188188 350593 193882 350829
rect 194118 350593 199813 350829
rect 200049 350593 215952 350829
rect 216188 350593 221882 350829
rect 222118 350593 227813 350829
rect 228049 350593 243952 350829
rect 244188 350593 249882 350829
rect 250118 350593 255813 350829
rect 256049 350593 271952 350829
rect 272188 350593 277882 350829
rect 278118 350593 283813 350829
rect 284049 350593 299952 350829
rect 300188 350593 305882 350829
rect 306118 350593 311813 350829
rect 312049 350593 327952 350829
rect 328188 350593 333882 350829
rect 334118 350593 339813 350829
rect 340049 350593 355952 350829
rect 356188 350593 361882 350829
rect 362118 350593 367813 350829
rect 368049 350593 383952 350829
rect 384188 350593 389882 350829
rect 390118 350593 395813 350829
rect 396049 350593 411952 350829
rect 412188 350593 417882 350829
rect 418118 350593 423813 350829
rect 424049 350593 439952 350829
rect 440188 350593 445882 350829
rect 446118 350593 451813 350829
rect 452049 350593 467952 350829
rect 468188 350593 473882 350829
rect 474118 350593 479813 350829
rect 480049 350593 495952 350829
rect 496188 350593 501882 350829
rect 502118 350593 507813 350829
rect 508049 350593 523952 350829
rect 524188 350593 529882 350829
rect 530118 350593 535813 350829
rect 536049 350593 551952 350829
rect 552188 350593 557882 350829
rect 558118 350593 563813 350829
rect 564049 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 592650 350829
rect -8726 350509 592650 350593
rect -8726 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 19952 350509
rect 20188 350273 25882 350509
rect 26118 350273 31813 350509
rect 32049 350273 47952 350509
rect 48188 350273 53882 350509
rect 54118 350273 59813 350509
rect 60049 350273 75952 350509
rect 76188 350273 81882 350509
rect 82118 350273 87813 350509
rect 88049 350273 103952 350509
rect 104188 350273 109882 350509
rect 110118 350273 115813 350509
rect 116049 350273 131952 350509
rect 132188 350273 137882 350509
rect 138118 350273 143813 350509
rect 144049 350273 159952 350509
rect 160188 350273 165882 350509
rect 166118 350273 171813 350509
rect 172049 350273 187952 350509
rect 188188 350273 193882 350509
rect 194118 350273 199813 350509
rect 200049 350273 215952 350509
rect 216188 350273 221882 350509
rect 222118 350273 227813 350509
rect 228049 350273 243952 350509
rect 244188 350273 249882 350509
rect 250118 350273 255813 350509
rect 256049 350273 271952 350509
rect 272188 350273 277882 350509
rect 278118 350273 283813 350509
rect 284049 350273 299952 350509
rect 300188 350273 305882 350509
rect 306118 350273 311813 350509
rect 312049 350273 327952 350509
rect 328188 350273 333882 350509
rect 334118 350273 339813 350509
rect 340049 350273 355952 350509
rect 356188 350273 361882 350509
rect 362118 350273 367813 350509
rect 368049 350273 383952 350509
rect 384188 350273 389882 350509
rect 390118 350273 395813 350509
rect 396049 350273 411952 350509
rect 412188 350273 417882 350509
rect 418118 350273 423813 350509
rect 424049 350273 439952 350509
rect 440188 350273 445882 350509
rect 446118 350273 451813 350509
rect 452049 350273 467952 350509
rect 468188 350273 473882 350509
rect 474118 350273 479813 350509
rect 480049 350273 495952 350509
rect 496188 350273 501882 350509
rect 502118 350273 507813 350509
rect 508049 350273 523952 350509
rect 524188 350273 529882 350509
rect 530118 350273 535813 350509
rect 536049 350273 551952 350509
rect 552188 350273 557882 350509
rect 558118 350273 563813 350509
rect 564049 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 592650 350509
rect -8726 350241 592650 350273
rect -8726 347454 592650 347486
rect -8726 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 22916 347454
rect 23152 347218 28847 347454
rect 29083 347218 50916 347454
rect 51152 347218 56847 347454
rect 57083 347218 78916 347454
rect 79152 347218 84847 347454
rect 85083 347218 106916 347454
rect 107152 347218 112847 347454
rect 113083 347218 134916 347454
rect 135152 347218 140847 347454
rect 141083 347218 162916 347454
rect 163152 347218 168847 347454
rect 169083 347218 190916 347454
rect 191152 347218 196847 347454
rect 197083 347218 218916 347454
rect 219152 347218 224847 347454
rect 225083 347218 246916 347454
rect 247152 347218 252847 347454
rect 253083 347218 274916 347454
rect 275152 347218 280847 347454
rect 281083 347218 302916 347454
rect 303152 347218 308847 347454
rect 309083 347218 330916 347454
rect 331152 347218 336847 347454
rect 337083 347218 358916 347454
rect 359152 347218 364847 347454
rect 365083 347218 386916 347454
rect 387152 347218 392847 347454
rect 393083 347218 414916 347454
rect 415152 347218 420847 347454
rect 421083 347218 442916 347454
rect 443152 347218 448847 347454
rect 449083 347218 470916 347454
rect 471152 347218 476847 347454
rect 477083 347218 498916 347454
rect 499152 347218 504847 347454
rect 505083 347218 526916 347454
rect 527152 347218 532847 347454
rect 533083 347218 554916 347454
rect 555152 347218 560847 347454
rect 561083 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 592650 347454
rect -8726 347134 592650 347218
rect -8726 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 22916 347134
rect 23152 346898 28847 347134
rect 29083 346898 50916 347134
rect 51152 346898 56847 347134
rect 57083 346898 78916 347134
rect 79152 346898 84847 347134
rect 85083 346898 106916 347134
rect 107152 346898 112847 347134
rect 113083 346898 134916 347134
rect 135152 346898 140847 347134
rect 141083 346898 162916 347134
rect 163152 346898 168847 347134
rect 169083 346898 190916 347134
rect 191152 346898 196847 347134
rect 197083 346898 218916 347134
rect 219152 346898 224847 347134
rect 225083 346898 246916 347134
rect 247152 346898 252847 347134
rect 253083 346898 274916 347134
rect 275152 346898 280847 347134
rect 281083 346898 302916 347134
rect 303152 346898 308847 347134
rect 309083 346898 330916 347134
rect 331152 346898 336847 347134
rect 337083 346898 358916 347134
rect 359152 346898 364847 347134
rect 365083 346898 386916 347134
rect 387152 346898 392847 347134
rect 393083 346898 414916 347134
rect 415152 346898 420847 347134
rect 421083 346898 442916 347134
rect 443152 346898 448847 347134
rect 449083 346898 470916 347134
rect 471152 346898 476847 347134
rect 477083 346898 498916 347134
rect 499152 346898 504847 347134
rect 505083 346898 526916 347134
rect 527152 346898 532847 347134
rect 533083 346898 554916 347134
rect 555152 346898 560847 347134
rect 561083 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 592650 347134
rect -8726 346866 592650 346898
rect -8726 323829 592650 323861
rect -8726 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 19952 323829
rect 20188 323593 25882 323829
rect 26118 323593 31813 323829
rect 32049 323593 47952 323829
rect 48188 323593 53882 323829
rect 54118 323593 59813 323829
rect 60049 323593 75952 323829
rect 76188 323593 81882 323829
rect 82118 323593 87813 323829
rect 88049 323593 103952 323829
rect 104188 323593 109882 323829
rect 110118 323593 115813 323829
rect 116049 323593 131952 323829
rect 132188 323593 137882 323829
rect 138118 323593 143813 323829
rect 144049 323593 159952 323829
rect 160188 323593 165882 323829
rect 166118 323593 171813 323829
rect 172049 323593 187952 323829
rect 188188 323593 193882 323829
rect 194118 323593 199813 323829
rect 200049 323593 215952 323829
rect 216188 323593 221882 323829
rect 222118 323593 227813 323829
rect 228049 323593 243952 323829
rect 244188 323593 249882 323829
rect 250118 323593 255813 323829
rect 256049 323593 271952 323829
rect 272188 323593 277882 323829
rect 278118 323593 283813 323829
rect 284049 323593 299952 323829
rect 300188 323593 305882 323829
rect 306118 323593 311813 323829
rect 312049 323593 327952 323829
rect 328188 323593 333882 323829
rect 334118 323593 339813 323829
rect 340049 323593 355952 323829
rect 356188 323593 361882 323829
rect 362118 323593 367813 323829
rect 368049 323593 383952 323829
rect 384188 323593 389882 323829
rect 390118 323593 395813 323829
rect 396049 323593 411952 323829
rect 412188 323593 417882 323829
rect 418118 323593 423813 323829
rect 424049 323593 439952 323829
rect 440188 323593 445882 323829
rect 446118 323593 451813 323829
rect 452049 323593 467952 323829
rect 468188 323593 473882 323829
rect 474118 323593 479813 323829
rect 480049 323593 495952 323829
rect 496188 323593 501882 323829
rect 502118 323593 507813 323829
rect 508049 323593 523952 323829
rect 524188 323593 529882 323829
rect 530118 323593 535813 323829
rect 536049 323593 551952 323829
rect 552188 323593 557882 323829
rect 558118 323593 563813 323829
rect 564049 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 592650 323829
rect -8726 323509 592650 323593
rect -8726 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 19952 323509
rect 20188 323273 25882 323509
rect 26118 323273 31813 323509
rect 32049 323273 47952 323509
rect 48188 323273 53882 323509
rect 54118 323273 59813 323509
rect 60049 323273 75952 323509
rect 76188 323273 81882 323509
rect 82118 323273 87813 323509
rect 88049 323273 103952 323509
rect 104188 323273 109882 323509
rect 110118 323273 115813 323509
rect 116049 323273 131952 323509
rect 132188 323273 137882 323509
rect 138118 323273 143813 323509
rect 144049 323273 159952 323509
rect 160188 323273 165882 323509
rect 166118 323273 171813 323509
rect 172049 323273 187952 323509
rect 188188 323273 193882 323509
rect 194118 323273 199813 323509
rect 200049 323273 215952 323509
rect 216188 323273 221882 323509
rect 222118 323273 227813 323509
rect 228049 323273 243952 323509
rect 244188 323273 249882 323509
rect 250118 323273 255813 323509
rect 256049 323273 271952 323509
rect 272188 323273 277882 323509
rect 278118 323273 283813 323509
rect 284049 323273 299952 323509
rect 300188 323273 305882 323509
rect 306118 323273 311813 323509
rect 312049 323273 327952 323509
rect 328188 323273 333882 323509
rect 334118 323273 339813 323509
rect 340049 323273 355952 323509
rect 356188 323273 361882 323509
rect 362118 323273 367813 323509
rect 368049 323273 383952 323509
rect 384188 323273 389882 323509
rect 390118 323273 395813 323509
rect 396049 323273 411952 323509
rect 412188 323273 417882 323509
rect 418118 323273 423813 323509
rect 424049 323273 439952 323509
rect 440188 323273 445882 323509
rect 446118 323273 451813 323509
rect 452049 323273 467952 323509
rect 468188 323273 473882 323509
rect 474118 323273 479813 323509
rect 480049 323273 495952 323509
rect 496188 323273 501882 323509
rect 502118 323273 507813 323509
rect 508049 323273 523952 323509
rect 524188 323273 529882 323509
rect 530118 323273 535813 323509
rect 536049 323273 551952 323509
rect 552188 323273 557882 323509
rect 558118 323273 563813 323509
rect 564049 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 592650 323509
rect -8726 323241 592650 323273
rect -8726 320454 592650 320486
rect -8726 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 22916 320454
rect 23152 320218 28847 320454
rect 29083 320218 50916 320454
rect 51152 320218 56847 320454
rect 57083 320218 78916 320454
rect 79152 320218 84847 320454
rect 85083 320218 106916 320454
rect 107152 320218 112847 320454
rect 113083 320218 134916 320454
rect 135152 320218 140847 320454
rect 141083 320218 162916 320454
rect 163152 320218 168847 320454
rect 169083 320218 190916 320454
rect 191152 320218 196847 320454
rect 197083 320218 218916 320454
rect 219152 320218 224847 320454
rect 225083 320218 246916 320454
rect 247152 320218 252847 320454
rect 253083 320218 274916 320454
rect 275152 320218 280847 320454
rect 281083 320218 302916 320454
rect 303152 320218 308847 320454
rect 309083 320218 330916 320454
rect 331152 320218 336847 320454
rect 337083 320218 358916 320454
rect 359152 320218 364847 320454
rect 365083 320218 386916 320454
rect 387152 320218 392847 320454
rect 393083 320218 414916 320454
rect 415152 320218 420847 320454
rect 421083 320218 442916 320454
rect 443152 320218 448847 320454
rect 449083 320218 470916 320454
rect 471152 320218 476847 320454
rect 477083 320218 498916 320454
rect 499152 320218 504847 320454
rect 505083 320218 526916 320454
rect 527152 320218 532847 320454
rect 533083 320218 554916 320454
rect 555152 320218 560847 320454
rect 561083 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 592650 320454
rect -8726 320134 592650 320218
rect -8726 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 22916 320134
rect 23152 319898 28847 320134
rect 29083 319898 50916 320134
rect 51152 319898 56847 320134
rect 57083 319898 78916 320134
rect 79152 319898 84847 320134
rect 85083 319898 106916 320134
rect 107152 319898 112847 320134
rect 113083 319898 134916 320134
rect 135152 319898 140847 320134
rect 141083 319898 162916 320134
rect 163152 319898 168847 320134
rect 169083 319898 190916 320134
rect 191152 319898 196847 320134
rect 197083 319898 218916 320134
rect 219152 319898 224847 320134
rect 225083 319898 246916 320134
rect 247152 319898 252847 320134
rect 253083 319898 274916 320134
rect 275152 319898 280847 320134
rect 281083 319898 302916 320134
rect 303152 319898 308847 320134
rect 309083 319898 330916 320134
rect 331152 319898 336847 320134
rect 337083 319898 358916 320134
rect 359152 319898 364847 320134
rect 365083 319898 386916 320134
rect 387152 319898 392847 320134
rect 393083 319898 414916 320134
rect 415152 319898 420847 320134
rect 421083 319898 442916 320134
rect 443152 319898 448847 320134
rect 449083 319898 470916 320134
rect 471152 319898 476847 320134
rect 477083 319898 498916 320134
rect 499152 319898 504847 320134
rect 505083 319898 526916 320134
rect 527152 319898 532847 320134
rect 533083 319898 554916 320134
rect 555152 319898 560847 320134
rect 561083 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 592650 320134
rect -8726 319866 592650 319898
rect -8726 296829 592650 296861
rect -8726 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 19952 296829
rect 20188 296593 25882 296829
rect 26118 296593 31813 296829
rect 32049 296593 47952 296829
rect 48188 296593 53882 296829
rect 54118 296593 59813 296829
rect 60049 296593 75952 296829
rect 76188 296593 81882 296829
rect 82118 296593 87813 296829
rect 88049 296593 103952 296829
rect 104188 296593 109882 296829
rect 110118 296593 115813 296829
rect 116049 296593 131952 296829
rect 132188 296593 137882 296829
rect 138118 296593 143813 296829
rect 144049 296593 159952 296829
rect 160188 296593 165882 296829
rect 166118 296593 171813 296829
rect 172049 296593 187952 296829
rect 188188 296593 193882 296829
rect 194118 296593 199813 296829
rect 200049 296593 215952 296829
rect 216188 296593 221882 296829
rect 222118 296593 227813 296829
rect 228049 296593 243952 296829
rect 244188 296593 249882 296829
rect 250118 296593 255813 296829
rect 256049 296593 271952 296829
rect 272188 296593 277882 296829
rect 278118 296593 283813 296829
rect 284049 296593 299952 296829
rect 300188 296593 305882 296829
rect 306118 296593 311813 296829
rect 312049 296593 327952 296829
rect 328188 296593 333882 296829
rect 334118 296593 339813 296829
rect 340049 296593 355952 296829
rect 356188 296593 361882 296829
rect 362118 296593 367813 296829
rect 368049 296593 383952 296829
rect 384188 296593 389882 296829
rect 390118 296593 395813 296829
rect 396049 296593 411952 296829
rect 412188 296593 417882 296829
rect 418118 296593 423813 296829
rect 424049 296593 439952 296829
rect 440188 296593 445882 296829
rect 446118 296593 451813 296829
rect 452049 296593 467952 296829
rect 468188 296593 473882 296829
rect 474118 296593 479813 296829
rect 480049 296593 495952 296829
rect 496188 296593 501882 296829
rect 502118 296593 507813 296829
rect 508049 296593 523952 296829
rect 524188 296593 529882 296829
rect 530118 296593 535813 296829
rect 536049 296593 551952 296829
rect 552188 296593 557882 296829
rect 558118 296593 563813 296829
rect 564049 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 592650 296829
rect -8726 296509 592650 296593
rect -8726 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 19952 296509
rect 20188 296273 25882 296509
rect 26118 296273 31813 296509
rect 32049 296273 47952 296509
rect 48188 296273 53882 296509
rect 54118 296273 59813 296509
rect 60049 296273 75952 296509
rect 76188 296273 81882 296509
rect 82118 296273 87813 296509
rect 88049 296273 103952 296509
rect 104188 296273 109882 296509
rect 110118 296273 115813 296509
rect 116049 296273 131952 296509
rect 132188 296273 137882 296509
rect 138118 296273 143813 296509
rect 144049 296273 159952 296509
rect 160188 296273 165882 296509
rect 166118 296273 171813 296509
rect 172049 296273 187952 296509
rect 188188 296273 193882 296509
rect 194118 296273 199813 296509
rect 200049 296273 215952 296509
rect 216188 296273 221882 296509
rect 222118 296273 227813 296509
rect 228049 296273 243952 296509
rect 244188 296273 249882 296509
rect 250118 296273 255813 296509
rect 256049 296273 271952 296509
rect 272188 296273 277882 296509
rect 278118 296273 283813 296509
rect 284049 296273 299952 296509
rect 300188 296273 305882 296509
rect 306118 296273 311813 296509
rect 312049 296273 327952 296509
rect 328188 296273 333882 296509
rect 334118 296273 339813 296509
rect 340049 296273 355952 296509
rect 356188 296273 361882 296509
rect 362118 296273 367813 296509
rect 368049 296273 383952 296509
rect 384188 296273 389882 296509
rect 390118 296273 395813 296509
rect 396049 296273 411952 296509
rect 412188 296273 417882 296509
rect 418118 296273 423813 296509
rect 424049 296273 439952 296509
rect 440188 296273 445882 296509
rect 446118 296273 451813 296509
rect 452049 296273 467952 296509
rect 468188 296273 473882 296509
rect 474118 296273 479813 296509
rect 480049 296273 495952 296509
rect 496188 296273 501882 296509
rect 502118 296273 507813 296509
rect 508049 296273 523952 296509
rect 524188 296273 529882 296509
rect 530118 296273 535813 296509
rect 536049 296273 551952 296509
rect 552188 296273 557882 296509
rect 558118 296273 563813 296509
rect 564049 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 592650 296509
rect -8726 296241 592650 296273
rect -8726 293454 592650 293486
rect -8726 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 22916 293454
rect 23152 293218 28847 293454
rect 29083 293218 50916 293454
rect 51152 293218 56847 293454
rect 57083 293218 78916 293454
rect 79152 293218 84847 293454
rect 85083 293218 106916 293454
rect 107152 293218 112847 293454
rect 113083 293218 134916 293454
rect 135152 293218 140847 293454
rect 141083 293218 162916 293454
rect 163152 293218 168847 293454
rect 169083 293218 190916 293454
rect 191152 293218 196847 293454
rect 197083 293218 218916 293454
rect 219152 293218 224847 293454
rect 225083 293218 246916 293454
rect 247152 293218 252847 293454
rect 253083 293218 274916 293454
rect 275152 293218 280847 293454
rect 281083 293218 302916 293454
rect 303152 293218 308847 293454
rect 309083 293218 330916 293454
rect 331152 293218 336847 293454
rect 337083 293218 358916 293454
rect 359152 293218 364847 293454
rect 365083 293218 386916 293454
rect 387152 293218 392847 293454
rect 393083 293218 414916 293454
rect 415152 293218 420847 293454
rect 421083 293218 442916 293454
rect 443152 293218 448847 293454
rect 449083 293218 470916 293454
rect 471152 293218 476847 293454
rect 477083 293218 498916 293454
rect 499152 293218 504847 293454
rect 505083 293218 526916 293454
rect 527152 293218 532847 293454
rect 533083 293218 554916 293454
rect 555152 293218 560847 293454
rect 561083 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 592650 293454
rect -8726 293134 592650 293218
rect -8726 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 22916 293134
rect 23152 292898 28847 293134
rect 29083 292898 50916 293134
rect 51152 292898 56847 293134
rect 57083 292898 78916 293134
rect 79152 292898 84847 293134
rect 85083 292898 106916 293134
rect 107152 292898 112847 293134
rect 113083 292898 134916 293134
rect 135152 292898 140847 293134
rect 141083 292898 162916 293134
rect 163152 292898 168847 293134
rect 169083 292898 190916 293134
rect 191152 292898 196847 293134
rect 197083 292898 218916 293134
rect 219152 292898 224847 293134
rect 225083 292898 246916 293134
rect 247152 292898 252847 293134
rect 253083 292898 274916 293134
rect 275152 292898 280847 293134
rect 281083 292898 302916 293134
rect 303152 292898 308847 293134
rect 309083 292898 330916 293134
rect 331152 292898 336847 293134
rect 337083 292898 358916 293134
rect 359152 292898 364847 293134
rect 365083 292898 386916 293134
rect 387152 292898 392847 293134
rect 393083 292898 414916 293134
rect 415152 292898 420847 293134
rect 421083 292898 442916 293134
rect 443152 292898 448847 293134
rect 449083 292898 470916 293134
rect 471152 292898 476847 293134
rect 477083 292898 498916 293134
rect 499152 292898 504847 293134
rect 505083 292898 526916 293134
rect 527152 292898 532847 293134
rect 533083 292898 554916 293134
rect 555152 292898 560847 293134
rect 561083 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 592650 293134
rect -8726 292866 592650 292898
rect -8726 269829 592650 269861
rect -8726 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 19952 269829
rect 20188 269593 25882 269829
rect 26118 269593 31813 269829
rect 32049 269593 47952 269829
rect 48188 269593 53882 269829
rect 54118 269593 59813 269829
rect 60049 269593 75952 269829
rect 76188 269593 81882 269829
rect 82118 269593 87813 269829
rect 88049 269593 103952 269829
rect 104188 269593 109882 269829
rect 110118 269593 115813 269829
rect 116049 269593 131952 269829
rect 132188 269593 137882 269829
rect 138118 269593 143813 269829
rect 144049 269593 159952 269829
rect 160188 269593 165882 269829
rect 166118 269593 171813 269829
rect 172049 269593 187952 269829
rect 188188 269593 193882 269829
rect 194118 269593 199813 269829
rect 200049 269593 215952 269829
rect 216188 269593 221882 269829
rect 222118 269593 227813 269829
rect 228049 269593 243952 269829
rect 244188 269593 249882 269829
rect 250118 269593 255813 269829
rect 256049 269593 271952 269829
rect 272188 269593 277882 269829
rect 278118 269593 283813 269829
rect 284049 269593 299952 269829
rect 300188 269593 305882 269829
rect 306118 269593 311813 269829
rect 312049 269593 327952 269829
rect 328188 269593 333882 269829
rect 334118 269593 339813 269829
rect 340049 269593 355952 269829
rect 356188 269593 361882 269829
rect 362118 269593 367813 269829
rect 368049 269593 383952 269829
rect 384188 269593 389882 269829
rect 390118 269593 395813 269829
rect 396049 269593 411952 269829
rect 412188 269593 417882 269829
rect 418118 269593 423813 269829
rect 424049 269593 439952 269829
rect 440188 269593 445882 269829
rect 446118 269593 451813 269829
rect 452049 269593 467952 269829
rect 468188 269593 473882 269829
rect 474118 269593 479813 269829
rect 480049 269593 495952 269829
rect 496188 269593 501882 269829
rect 502118 269593 507813 269829
rect 508049 269593 523952 269829
rect 524188 269593 529882 269829
rect 530118 269593 535813 269829
rect 536049 269593 551952 269829
rect 552188 269593 557882 269829
rect 558118 269593 563813 269829
rect 564049 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 592650 269829
rect -8726 269509 592650 269593
rect -8726 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 19952 269509
rect 20188 269273 25882 269509
rect 26118 269273 31813 269509
rect 32049 269273 47952 269509
rect 48188 269273 53882 269509
rect 54118 269273 59813 269509
rect 60049 269273 75952 269509
rect 76188 269273 81882 269509
rect 82118 269273 87813 269509
rect 88049 269273 103952 269509
rect 104188 269273 109882 269509
rect 110118 269273 115813 269509
rect 116049 269273 131952 269509
rect 132188 269273 137882 269509
rect 138118 269273 143813 269509
rect 144049 269273 159952 269509
rect 160188 269273 165882 269509
rect 166118 269273 171813 269509
rect 172049 269273 187952 269509
rect 188188 269273 193882 269509
rect 194118 269273 199813 269509
rect 200049 269273 215952 269509
rect 216188 269273 221882 269509
rect 222118 269273 227813 269509
rect 228049 269273 243952 269509
rect 244188 269273 249882 269509
rect 250118 269273 255813 269509
rect 256049 269273 271952 269509
rect 272188 269273 277882 269509
rect 278118 269273 283813 269509
rect 284049 269273 299952 269509
rect 300188 269273 305882 269509
rect 306118 269273 311813 269509
rect 312049 269273 327952 269509
rect 328188 269273 333882 269509
rect 334118 269273 339813 269509
rect 340049 269273 355952 269509
rect 356188 269273 361882 269509
rect 362118 269273 367813 269509
rect 368049 269273 383952 269509
rect 384188 269273 389882 269509
rect 390118 269273 395813 269509
rect 396049 269273 411952 269509
rect 412188 269273 417882 269509
rect 418118 269273 423813 269509
rect 424049 269273 439952 269509
rect 440188 269273 445882 269509
rect 446118 269273 451813 269509
rect 452049 269273 467952 269509
rect 468188 269273 473882 269509
rect 474118 269273 479813 269509
rect 480049 269273 495952 269509
rect 496188 269273 501882 269509
rect 502118 269273 507813 269509
rect 508049 269273 523952 269509
rect 524188 269273 529882 269509
rect 530118 269273 535813 269509
rect 536049 269273 551952 269509
rect 552188 269273 557882 269509
rect 558118 269273 563813 269509
rect 564049 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 592650 269509
rect -8726 269241 592650 269273
rect -8726 266454 592650 266486
rect -8726 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 22916 266454
rect 23152 266218 28847 266454
rect 29083 266218 50916 266454
rect 51152 266218 56847 266454
rect 57083 266218 78916 266454
rect 79152 266218 84847 266454
rect 85083 266218 106916 266454
rect 107152 266218 112847 266454
rect 113083 266218 134916 266454
rect 135152 266218 140847 266454
rect 141083 266218 162916 266454
rect 163152 266218 168847 266454
rect 169083 266218 190916 266454
rect 191152 266218 196847 266454
rect 197083 266218 218916 266454
rect 219152 266218 224847 266454
rect 225083 266218 246916 266454
rect 247152 266218 252847 266454
rect 253083 266218 274916 266454
rect 275152 266218 280847 266454
rect 281083 266218 302916 266454
rect 303152 266218 308847 266454
rect 309083 266218 330916 266454
rect 331152 266218 336847 266454
rect 337083 266218 358916 266454
rect 359152 266218 364847 266454
rect 365083 266218 386916 266454
rect 387152 266218 392847 266454
rect 393083 266218 414916 266454
rect 415152 266218 420847 266454
rect 421083 266218 442916 266454
rect 443152 266218 448847 266454
rect 449083 266218 470916 266454
rect 471152 266218 476847 266454
rect 477083 266218 498916 266454
rect 499152 266218 504847 266454
rect 505083 266218 526916 266454
rect 527152 266218 532847 266454
rect 533083 266218 554916 266454
rect 555152 266218 560847 266454
rect 561083 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 592650 266454
rect -8726 266134 592650 266218
rect -8726 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 22916 266134
rect 23152 265898 28847 266134
rect 29083 265898 50916 266134
rect 51152 265898 56847 266134
rect 57083 265898 78916 266134
rect 79152 265898 84847 266134
rect 85083 265898 106916 266134
rect 107152 265898 112847 266134
rect 113083 265898 134916 266134
rect 135152 265898 140847 266134
rect 141083 265898 162916 266134
rect 163152 265898 168847 266134
rect 169083 265898 190916 266134
rect 191152 265898 196847 266134
rect 197083 265898 218916 266134
rect 219152 265898 224847 266134
rect 225083 265898 246916 266134
rect 247152 265898 252847 266134
rect 253083 265898 274916 266134
rect 275152 265898 280847 266134
rect 281083 265898 302916 266134
rect 303152 265898 308847 266134
rect 309083 265898 330916 266134
rect 331152 265898 336847 266134
rect 337083 265898 358916 266134
rect 359152 265898 364847 266134
rect 365083 265898 386916 266134
rect 387152 265898 392847 266134
rect 393083 265898 414916 266134
rect 415152 265898 420847 266134
rect 421083 265898 442916 266134
rect 443152 265898 448847 266134
rect 449083 265898 470916 266134
rect 471152 265898 476847 266134
rect 477083 265898 498916 266134
rect 499152 265898 504847 266134
rect 505083 265898 526916 266134
rect 527152 265898 532847 266134
rect 533083 265898 554916 266134
rect 555152 265898 560847 266134
rect 561083 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 592650 266134
rect -8726 265866 592650 265898
rect -8726 242829 592650 242861
rect -8726 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 19952 242829
rect 20188 242593 25882 242829
rect 26118 242593 31813 242829
rect 32049 242593 47952 242829
rect 48188 242593 53882 242829
rect 54118 242593 59813 242829
rect 60049 242593 75952 242829
rect 76188 242593 81882 242829
rect 82118 242593 87813 242829
rect 88049 242593 103952 242829
rect 104188 242593 109882 242829
rect 110118 242593 115813 242829
rect 116049 242593 131952 242829
rect 132188 242593 137882 242829
rect 138118 242593 143813 242829
rect 144049 242593 159952 242829
rect 160188 242593 165882 242829
rect 166118 242593 171813 242829
rect 172049 242593 187952 242829
rect 188188 242593 193882 242829
rect 194118 242593 199813 242829
rect 200049 242593 215952 242829
rect 216188 242593 221882 242829
rect 222118 242593 227813 242829
rect 228049 242593 243952 242829
rect 244188 242593 249882 242829
rect 250118 242593 255813 242829
rect 256049 242593 271952 242829
rect 272188 242593 277882 242829
rect 278118 242593 283813 242829
rect 284049 242593 299952 242829
rect 300188 242593 305882 242829
rect 306118 242593 311813 242829
rect 312049 242593 327952 242829
rect 328188 242593 333882 242829
rect 334118 242593 339813 242829
rect 340049 242593 355952 242829
rect 356188 242593 361882 242829
rect 362118 242593 367813 242829
rect 368049 242593 383952 242829
rect 384188 242593 389882 242829
rect 390118 242593 395813 242829
rect 396049 242593 411952 242829
rect 412188 242593 417882 242829
rect 418118 242593 423813 242829
rect 424049 242593 439952 242829
rect 440188 242593 445882 242829
rect 446118 242593 451813 242829
rect 452049 242593 467952 242829
rect 468188 242593 473882 242829
rect 474118 242593 479813 242829
rect 480049 242593 495952 242829
rect 496188 242593 501882 242829
rect 502118 242593 507813 242829
rect 508049 242593 523952 242829
rect 524188 242593 529882 242829
rect 530118 242593 535813 242829
rect 536049 242593 551952 242829
rect 552188 242593 557882 242829
rect 558118 242593 563813 242829
rect 564049 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 592650 242829
rect -8726 242509 592650 242593
rect -8726 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 19952 242509
rect 20188 242273 25882 242509
rect 26118 242273 31813 242509
rect 32049 242273 47952 242509
rect 48188 242273 53882 242509
rect 54118 242273 59813 242509
rect 60049 242273 75952 242509
rect 76188 242273 81882 242509
rect 82118 242273 87813 242509
rect 88049 242273 103952 242509
rect 104188 242273 109882 242509
rect 110118 242273 115813 242509
rect 116049 242273 131952 242509
rect 132188 242273 137882 242509
rect 138118 242273 143813 242509
rect 144049 242273 159952 242509
rect 160188 242273 165882 242509
rect 166118 242273 171813 242509
rect 172049 242273 187952 242509
rect 188188 242273 193882 242509
rect 194118 242273 199813 242509
rect 200049 242273 215952 242509
rect 216188 242273 221882 242509
rect 222118 242273 227813 242509
rect 228049 242273 243952 242509
rect 244188 242273 249882 242509
rect 250118 242273 255813 242509
rect 256049 242273 271952 242509
rect 272188 242273 277882 242509
rect 278118 242273 283813 242509
rect 284049 242273 299952 242509
rect 300188 242273 305882 242509
rect 306118 242273 311813 242509
rect 312049 242273 327952 242509
rect 328188 242273 333882 242509
rect 334118 242273 339813 242509
rect 340049 242273 355952 242509
rect 356188 242273 361882 242509
rect 362118 242273 367813 242509
rect 368049 242273 383952 242509
rect 384188 242273 389882 242509
rect 390118 242273 395813 242509
rect 396049 242273 411952 242509
rect 412188 242273 417882 242509
rect 418118 242273 423813 242509
rect 424049 242273 439952 242509
rect 440188 242273 445882 242509
rect 446118 242273 451813 242509
rect 452049 242273 467952 242509
rect 468188 242273 473882 242509
rect 474118 242273 479813 242509
rect 480049 242273 495952 242509
rect 496188 242273 501882 242509
rect 502118 242273 507813 242509
rect 508049 242273 523952 242509
rect 524188 242273 529882 242509
rect 530118 242273 535813 242509
rect 536049 242273 551952 242509
rect 552188 242273 557882 242509
rect 558118 242273 563813 242509
rect 564049 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 592650 242509
rect -8726 242241 592650 242273
rect -8726 239454 592650 239486
rect -8726 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 22916 239454
rect 23152 239218 28847 239454
rect 29083 239218 50916 239454
rect 51152 239218 56847 239454
rect 57083 239218 78916 239454
rect 79152 239218 84847 239454
rect 85083 239218 106916 239454
rect 107152 239218 112847 239454
rect 113083 239218 134916 239454
rect 135152 239218 140847 239454
rect 141083 239218 162916 239454
rect 163152 239218 168847 239454
rect 169083 239218 190916 239454
rect 191152 239218 196847 239454
rect 197083 239218 218916 239454
rect 219152 239218 224847 239454
rect 225083 239218 246916 239454
rect 247152 239218 252847 239454
rect 253083 239218 274916 239454
rect 275152 239218 280847 239454
rect 281083 239218 302916 239454
rect 303152 239218 308847 239454
rect 309083 239218 330916 239454
rect 331152 239218 336847 239454
rect 337083 239218 358916 239454
rect 359152 239218 364847 239454
rect 365083 239218 386916 239454
rect 387152 239218 392847 239454
rect 393083 239218 414916 239454
rect 415152 239218 420847 239454
rect 421083 239218 442916 239454
rect 443152 239218 448847 239454
rect 449083 239218 470916 239454
rect 471152 239218 476847 239454
rect 477083 239218 498916 239454
rect 499152 239218 504847 239454
rect 505083 239218 526916 239454
rect 527152 239218 532847 239454
rect 533083 239218 554916 239454
rect 555152 239218 560847 239454
rect 561083 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 592650 239454
rect -8726 239134 592650 239218
rect -8726 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 22916 239134
rect 23152 238898 28847 239134
rect 29083 238898 50916 239134
rect 51152 238898 56847 239134
rect 57083 238898 78916 239134
rect 79152 238898 84847 239134
rect 85083 238898 106916 239134
rect 107152 238898 112847 239134
rect 113083 238898 134916 239134
rect 135152 238898 140847 239134
rect 141083 238898 162916 239134
rect 163152 238898 168847 239134
rect 169083 238898 190916 239134
rect 191152 238898 196847 239134
rect 197083 238898 218916 239134
rect 219152 238898 224847 239134
rect 225083 238898 246916 239134
rect 247152 238898 252847 239134
rect 253083 238898 274916 239134
rect 275152 238898 280847 239134
rect 281083 238898 302916 239134
rect 303152 238898 308847 239134
rect 309083 238898 330916 239134
rect 331152 238898 336847 239134
rect 337083 238898 358916 239134
rect 359152 238898 364847 239134
rect 365083 238898 386916 239134
rect 387152 238898 392847 239134
rect 393083 238898 414916 239134
rect 415152 238898 420847 239134
rect 421083 238898 442916 239134
rect 443152 238898 448847 239134
rect 449083 238898 470916 239134
rect 471152 238898 476847 239134
rect 477083 238898 498916 239134
rect 499152 238898 504847 239134
rect 505083 238898 526916 239134
rect 527152 238898 532847 239134
rect 533083 238898 554916 239134
rect 555152 238898 560847 239134
rect 561083 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 592650 239134
rect -8726 238866 592650 238898
rect -8726 215829 592650 215861
rect -8726 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 19952 215829
rect 20188 215593 25882 215829
rect 26118 215593 31813 215829
rect 32049 215593 47952 215829
rect 48188 215593 53882 215829
rect 54118 215593 59813 215829
rect 60049 215593 75952 215829
rect 76188 215593 81882 215829
rect 82118 215593 87813 215829
rect 88049 215593 103952 215829
rect 104188 215593 109882 215829
rect 110118 215593 115813 215829
rect 116049 215593 131952 215829
rect 132188 215593 137882 215829
rect 138118 215593 143813 215829
rect 144049 215593 159952 215829
rect 160188 215593 165882 215829
rect 166118 215593 171813 215829
rect 172049 215593 187952 215829
rect 188188 215593 193882 215829
rect 194118 215593 199813 215829
rect 200049 215593 215952 215829
rect 216188 215593 221882 215829
rect 222118 215593 227813 215829
rect 228049 215593 243952 215829
rect 244188 215593 249882 215829
rect 250118 215593 255813 215829
rect 256049 215593 271952 215829
rect 272188 215593 277882 215829
rect 278118 215593 283813 215829
rect 284049 215593 299952 215829
rect 300188 215593 305882 215829
rect 306118 215593 311813 215829
rect 312049 215593 327952 215829
rect 328188 215593 333882 215829
rect 334118 215593 339813 215829
rect 340049 215593 355952 215829
rect 356188 215593 361882 215829
rect 362118 215593 367813 215829
rect 368049 215593 383952 215829
rect 384188 215593 389882 215829
rect 390118 215593 395813 215829
rect 396049 215593 411952 215829
rect 412188 215593 417882 215829
rect 418118 215593 423813 215829
rect 424049 215593 439952 215829
rect 440188 215593 445882 215829
rect 446118 215593 451813 215829
rect 452049 215593 467952 215829
rect 468188 215593 473882 215829
rect 474118 215593 479813 215829
rect 480049 215593 495952 215829
rect 496188 215593 501882 215829
rect 502118 215593 507813 215829
rect 508049 215593 523952 215829
rect 524188 215593 529882 215829
rect 530118 215593 535813 215829
rect 536049 215593 551952 215829
rect 552188 215593 557882 215829
rect 558118 215593 563813 215829
rect 564049 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 592650 215829
rect -8726 215509 592650 215593
rect -8726 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 19952 215509
rect 20188 215273 25882 215509
rect 26118 215273 31813 215509
rect 32049 215273 47952 215509
rect 48188 215273 53882 215509
rect 54118 215273 59813 215509
rect 60049 215273 75952 215509
rect 76188 215273 81882 215509
rect 82118 215273 87813 215509
rect 88049 215273 103952 215509
rect 104188 215273 109882 215509
rect 110118 215273 115813 215509
rect 116049 215273 131952 215509
rect 132188 215273 137882 215509
rect 138118 215273 143813 215509
rect 144049 215273 159952 215509
rect 160188 215273 165882 215509
rect 166118 215273 171813 215509
rect 172049 215273 187952 215509
rect 188188 215273 193882 215509
rect 194118 215273 199813 215509
rect 200049 215273 215952 215509
rect 216188 215273 221882 215509
rect 222118 215273 227813 215509
rect 228049 215273 243952 215509
rect 244188 215273 249882 215509
rect 250118 215273 255813 215509
rect 256049 215273 271952 215509
rect 272188 215273 277882 215509
rect 278118 215273 283813 215509
rect 284049 215273 299952 215509
rect 300188 215273 305882 215509
rect 306118 215273 311813 215509
rect 312049 215273 327952 215509
rect 328188 215273 333882 215509
rect 334118 215273 339813 215509
rect 340049 215273 355952 215509
rect 356188 215273 361882 215509
rect 362118 215273 367813 215509
rect 368049 215273 383952 215509
rect 384188 215273 389882 215509
rect 390118 215273 395813 215509
rect 396049 215273 411952 215509
rect 412188 215273 417882 215509
rect 418118 215273 423813 215509
rect 424049 215273 439952 215509
rect 440188 215273 445882 215509
rect 446118 215273 451813 215509
rect 452049 215273 467952 215509
rect 468188 215273 473882 215509
rect 474118 215273 479813 215509
rect 480049 215273 495952 215509
rect 496188 215273 501882 215509
rect 502118 215273 507813 215509
rect 508049 215273 523952 215509
rect 524188 215273 529882 215509
rect 530118 215273 535813 215509
rect 536049 215273 551952 215509
rect 552188 215273 557882 215509
rect 558118 215273 563813 215509
rect 564049 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 592650 215509
rect -8726 215241 592650 215273
rect -8726 212454 592650 212486
rect -8726 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 22916 212454
rect 23152 212218 28847 212454
rect 29083 212218 50916 212454
rect 51152 212218 56847 212454
rect 57083 212218 78916 212454
rect 79152 212218 84847 212454
rect 85083 212218 106916 212454
rect 107152 212218 112847 212454
rect 113083 212218 134916 212454
rect 135152 212218 140847 212454
rect 141083 212218 162916 212454
rect 163152 212218 168847 212454
rect 169083 212218 190916 212454
rect 191152 212218 196847 212454
rect 197083 212218 218916 212454
rect 219152 212218 224847 212454
rect 225083 212218 246916 212454
rect 247152 212218 252847 212454
rect 253083 212218 274916 212454
rect 275152 212218 280847 212454
rect 281083 212218 302916 212454
rect 303152 212218 308847 212454
rect 309083 212218 330916 212454
rect 331152 212218 336847 212454
rect 337083 212218 358916 212454
rect 359152 212218 364847 212454
rect 365083 212218 386916 212454
rect 387152 212218 392847 212454
rect 393083 212218 414916 212454
rect 415152 212218 420847 212454
rect 421083 212218 442916 212454
rect 443152 212218 448847 212454
rect 449083 212218 470916 212454
rect 471152 212218 476847 212454
rect 477083 212218 498916 212454
rect 499152 212218 504847 212454
rect 505083 212218 526916 212454
rect 527152 212218 532847 212454
rect 533083 212218 554916 212454
rect 555152 212218 560847 212454
rect 561083 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 592650 212454
rect -8726 212134 592650 212218
rect -8726 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 22916 212134
rect 23152 211898 28847 212134
rect 29083 211898 50916 212134
rect 51152 211898 56847 212134
rect 57083 211898 78916 212134
rect 79152 211898 84847 212134
rect 85083 211898 106916 212134
rect 107152 211898 112847 212134
rect 113083 211898 134916 212134
rect 135152 211898 140847 212134
rect 141083 211898 162916 212134
rect 163152 211898 168847 212134
rect 169083 211898 190916 212134
rect 191152 211898 196847 212134
rect 197083 211898 218916 212134
rect 219152 211898 224847 212134
rect 225083 211898 246916 212134
rect 247152 211898 252847 212134
rect 253083 211898 274916 212134
rect 275152 211898 280847 212134
rect 281083 211898 302916 212134
rect 303152 211898 308847 212134
rect 309083 211898 330916 212134
rect 331152 211898 336847 212134
rect 337083 211898 358916 212134
rect 359152 211898 364847 212134
rect 365083 211898 386916 212134
rect 387152 211898 392847 212134
rect 393083 211898 414916 212134
rect 415152 211898 420847 212134
rect 421083 211898 442916 212134
rect 443152 211898 448847 212134
rect 449083 211898 470916 212134
rect 471152 211898 476847 212134
rect 477083 211898 498916 212134
rect 499152 211898 504847 212134
rect 505083 211898 526916 212134
rect 527152 211898 532847 212134
rect 533083 211898 554916 212134
rect 555152 211898 560847 212134
rect 561083 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 592650 212134
rect -8726 211866 592650 211898
rect -8726 188829 592650 188861
rect -8726 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 19952 188829
rect 20188 188593 25882 188829
rect 26118 188593 31813 188829
rect 32049 188593 47952 188829
rect 48188 188593 53882 188829
rect 54118 188593 59813 188829
rect 60049 188593 75952 188829
rect 76188 188593 81882 188829
rect 82118 188593 87813 188829
rect 88049 188593 103952 188829
rect 104188 188593 109882 188829
rect 110118 188593 115813 188829
rect 116049 188593 131952 188829
rect 132188 188593 137882 188829
rect 138118 188593 143813 188829
rect 144049 188593 159952 188829
rect 160188 188593 165882 188829
rect 166118 188593 171813 188829
rect 172049 188593 187952 188829
rect 188188 188593 193882 188829
rect 194118 188593 199813 188829
rect 200049 188593 215952 188829
rect 216188 188593 221882 188829
rect 222118 188593 227813 188829
rect 228049 188593 243952 188829
rect 244188 188593 249882 188829
rect 250118 188593 255813 188829
rect 256049 188593 271952 188829
rect 272188 188593 277882 188829
rect 278118 188593 283813 188829
rect 284049 188593 299952 188829
rect 300188 188593 305882 188829
rect 306118 188593 311813 188829
rect 312049 188593 327952 188829
rect 328188 188593 333882 188829
rect 334118 188593 339813 188829
rect 340049 188593 355952 188829
rect 356188 188593 361882 188829
rect 362118 188593 367813 188829
rect 368049 188593 383952 188829
rect 384188 188593 389882 188829
rect 390118 188593 395813 188829
rect 396049 188593 411952 188829
rect 412188 188593 417882 188829
rect 418118 188593 423813 188829
rect 424049 188593 439952 188829
rect 440188 188593 445882 188829
rect 446118 188593 451813 188829
rect 452049 188593 467952 188829
rect 468188 188593 473882 188829
rect 474118 188593 479813 188829
rect 480049 188593 495952 188829
rect 496188 188593 501882 188829
rect 502118 188593 507813 188829
rect 508049 188593 523952 188829
rect 524188 188593 529882 188829
rect 530118 188593 535813 188829
rect 536049 188593 551952 188829
rect 552188 188593 557882 188829
rect 558118 188593 563813 188829
rect 564049 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 592650 188829
rect -8726 188509 592650 188593
rect -8726 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 19952 188509
rect 20188 188273 25882 188509
rect 26118 188273 31813 188509
rect 32049 188273 47952 188509
rect 48188 188273 53882 188509
rect 54118 188273 59813 188509
rect 60049 188273 75952 188509
rect 76188 188273 81882 188509
rect 82118 188273 87813 188509
rect 88049 188273 103952 188509
rect 104188 188273 109882 188509
rect 110118 188273 115813 188509
rect 116049 188273 131952 188509
rect 132188 188273 137882 188509
rect 138118 188273 143813 188509
rect 144049 188273 159952 188509
rect 160188 188273 165882 188509
rect 166118 188273 171813 188509
rect 172049 188273 187952 188509
rect 188188 188273 193882 188509
rect 194118 188273 199813 188509
rect 200049 188273 215952 188509
rect 216188 188273 221882 188509
rect 222118 188273 227813 188509
rect 228049 188273 243952 188509
rect 244188 188273 249882 188509
rect 250118 188273 255813 188509
rect 256049 188273 271952 188509
rect 272188 188273 277882 188509
rect 278118 188273 283813 188509
rect 284049 188273 299952 188509
rect 300188 188273 305882 188509
rect 306118 188273 311813 188509
rect 312049 188273 327952 188509
rect 328188 188273 333882 188509
rect 334118 188273 339813 188509
rect 340049 188273 355952 188509
rect 356188 188273 361882 188509
rect 362118 188273 367813 188509
rect 368049 188273 383952 188509
rect 384188 188273 389882 188509
rect 390118 188273 395813 188509
rect 396049 188273 411952 188509
rect 412188 188273 417882 188509
rect 418118 188273 423813 188509
rect 424049 188273 439952 188509
rect 440188 188273 445882 188509
rect 446118 188273 451813 188509
rect 452049 188273 467952 188509
rect 468188 188273 473882 188509
rect 474118 188273 479813 188509
rect 480049 188273 495952 188509
rect 496188 188273 501882 188509
rect 502118 188273 507813 188509
rect 508049 188273 523952 188509
rect 524188 188273 529882 188509
rect 530118 188273 535813 188509
rect 536049 188273 551952 188509
rect 552188 188273 557882 188509
rect 558118 188273 563813 188509
rect 564049 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 592650 188509
rect -8726 188241 592650 188273
rect -8726 185454 592650 185486
rect -8726 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 22916 185454
rect 23152 185218 28847 185454
rect 29083 185218 50916 185454
rect 51152 185218 56847 185454
rect 57083 185218 78916 185454
rect 79152 185218 84847 185454
rect 85083 185218 106916 185454
rect 107152 185218 112847 185454
rect 113083 185218 134916 185454
rect 135152 185218 140847 185454
rect 141083 185218 162916 185454
rect 163152 185218 168847 185454
rect 169083 185218 190916 185454
rect 191152 185218 196847 185454
rect 197083 185218 218916 185454
rect 219152 185218 224847 185454
rect 225083 185218 246916 185454
rect 247152 185218 252847 185454
rect 253083 185218 274916 185454
rect 275152 185218 280847 185454
rect 281083 185218 302916 185454
rect 303152 185218 308847 185454
rect 309083 185218 330916 185454
rect 331152 185218 336847 185454
rect 337083 185218 358916 185454
rect 359152 185218 364847 185454
rect 365083 185218 386916 185454
rect 387152 185218 392847 185454
rect 393083 185218 414916 185454
rect 415152 185218 420847 185454
rect 421083 185218 442916 185454
rect 443152 185218 448847 185454
rect 449083 185218 470916 185454
rect 471152 185218 476847 185454
rect 477083 185218 498916 185454
rect 499152 185218 504847 185454
rect 505083 185218 526916 185454
rect 527152 185218 532847 185454
rect 533083 185218 554916 185454
rect 555152 185218 560847 185454
rect 561083 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 592650 185454
rect -8726 185134 592650 185218
rect -8726 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 22916 185134
rect 23152 184898 28847 185134
rect 29083 184898 50916 185134
rect 51152 184898 56847 185134
rect 57083 184898 78916 185134
rect 79152 184898 84847 185134
rect 85083 184898 106916 185134
rect 107152 184898 112847 185134
rect 113083 184898 134916 185134
rect 135152 184898 140847 185134
rect 141083 184898 162916 185134
rect 163152 184898 168847 185134
rect 169083 184898 190916 185134
rect 191152 184898 196847 185134
rect 197083 184898 218916 185134
rect 219152 184898 224847 185134
rect 225083 184898 246916 185134
rect 247152 184898 252847 185134
rect 253083 184898 274916 185134
rect 275152 184898 280847 185134
rect 281083 184898 302916 185134
rect 303152 184898 308847 185134
rect 309083 184898 330916 185134
rect 331152 184898 336847 185134
rect 337083 184898 358916 185134
rect 359152 184898 364847 185134
rect 365083 184898 386916 185134
rect 387152 184898 392847 185134
rect 393083 184898 414916 185134
rect 415152 184898 420847 185134
rect 421083 184898 442916 185134
rect 443152 184898 448847 185134
rect 449083 184898 470916 185134
rect 471152 184898 476847 185134
rect 477083 184898 498916 185134
rect 499152 184898 504847 185134
rect 505083 184898 526916 185134
rect 527152 184898 532847 185134
rect 533083 184898 554916 185134
rect 555152 184898 560847 185134
rect 561083 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 592650 185134
rect -8726 184866 592650 184898
rect -8726 161829 592650 161861
rect -8726 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 19952 161829
rect 20188 161593 25882 161829
rect 26118 161593 31813 161829
rect 32049 161593 47952 161829
rect 48188 161593 53882 161829
rect 54118 161593 59813 161829
rect 60049 161593 75952 161829
rect 76188 161593 81882 161829
rect 82118 161593 87813 161829
rect 88049 161593 103952 161829
rect 104188 161593 109882 161829
rect 110118 161593 115813 161829
rect 116049 161593 131952 161829
rect 132188 161593 137882 161829
rect 138118 161593 143813 161829
rect 144049 161593 159952 161829
rect 160188 161593 165882 161829
rect 166118 161593 171813 161829
rect 172049 161593 187952 161829
rect 188188 161593 193882 161829
rect 194118 161593 199813 161829
rect 200049 161593 215952 161829
rect 216188 161593 221882 161829
rect 222118 161593 227813 161829
rect 228049 161593 243952 161829
rect 244188 161593 249882 161829
rect 250118 161593 255813 161829
rect 256049 161593 271952 161829
rect 272188 161593 277882 161829
rect 278118 161593 283813 161829
rect 284049 161593 299952 161829
rect 300188 161593 305882 161829
rect 306118 161593 311813 161829
rect 312049 161593 327952 161829
rect 328188 161593 333882 161829
rect 334118 161593 339813 161829
rect 340049 161593 355952 161829
rect 356188 161593 361882 161829
rect 362118 161593 367813 161829
rect 368049 161593 383952 161829
rect 384188 161593 389882 161829
rect 390118 161593 395813 161829
rect 396049 161593 411952 161829
rect 412188 161593 417882 161829
rect 418118 161593 423813 161829
rect 424049 161593 439952 161829
rect 440188 161593 445882 161829
rect 446118 161593 451813 161829
rect 452049 161593 467952 161829
rect 468188 161593 473882 161829
rect 474118 161593 479813 161829
rect 480049 161593 495952 161829
rect 496188 161593 501882 161829
rect 502118 161593 507813 161829
rect 508049 161593 523952 161829
rect 524188 161593 529882 161829
rect 530118 161593 535813 161829
rect 536049 161593 551952 161829
rect 552188 161593 557882 161829
rect 558118 161593 563813 161829
rect 564049 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 592650 161829
rect -8726 161509 592650 161593
rect -8726 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 19952 161509
rect 20188 161273 25882 161509
rect 26118 161273 31813 161509
rect 32049 161273 47952 161509
rect 48188 161273 53882 161509
rect 54118 161273 59813 161509
rect 60049 161273 75952 161509
rect 76188 161273 81882 161509
rect 82118 161273 87813 161509
rect 88049 161273 103952 161509
rect 104188 161273 109882 161509
rect 110118 161273 115813 161509
rect 116049 161273 131952 161509
rect 132188 161273 137882 161509
rect 138118 161273 143813 161509
rect 144049 161273 159952 161509
rect 160188 161273 165882 161509
rect 166118 161273 171813 161509
rect 172049 161273 187952 161509
rect 188188 161273 193882 161509
rect 194118 161273 199813 161509
rect 200049 161273 215952 161509
rect 216188 161273 221882 161509
rect 222118 161273 227813 161509
rect 228049 161273 243952 161509
rect 244188 161273 249882 161509
rect 250118 161273 255813 161509
rect 256049 161273 271952 161509
rect 272188 161273 277882 161509
rect 278118 161273 283813 161509
rect 284049 161273 299952 161509
rect 300188 161273 305882 161509
rect 306118 161273 311813 161509
rect 312049 161273 327952 161509
rect 328188 161273 333882 161509
rect 334118 161273 339813 161509
rect 340049 161273 355952 161509
rect 356188 161273 361882 161509
rect 362118 161273 367813 161509
rect 368049 161273 383952 161509
rect 384188 161273 389882 161509
rect 390118 161273 395813 161509
rect 396049 161273 411952 161509
rect 412188 161273 417882 161509
rect 418118 161273 423813 161509
rect 424049 161273 439952 161509
rect 440188 161273 445882 161509
rect 446118 161273 451813 161509
rect 452049 161273 467952 161509
rect 468188 161273 473882 161509
rect 474118 161273 479813 161509
rect 480049 161273 495952 161509
rect 496188 161273 501882 161509
rect 502118 161273 507813 161509
rect 508049 161273 523952 161509
rect 524188 161273 529882 161509
rect 530118 161273 535813 161509
rect 536049 161273 551952 161509
rect 552188 161273 557882 161509
rect 558118 161273 563813 161509
rect 564049 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 592650 161509
rect -8726 161241 592650 161273
rect -8726 158454 592650 158486
rect -8726 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 22916 158454
rect 23152 158218 28847 158454
rect 29083 158218 50916 158454
rect 51152 158218 56847 158454
rect 57083 158218 78916 158454
rect 79152 158218 84847 158454
rect 85083 158218 106916 158454
rect 107152 158218 112847 158454
rect 113083 158218 134916 158454
rect 135152 158218 140847 158454
rect 141083 158218 162916 158454
rect 163152 158218 168847 158454
rect 169083 158218 190916 158454
rect 191152 158218 196847 158454
rect 197083 158218 218916 158454
rect 219152 158218 224847 158454
rect 225083 158218 246916 158454
rect 247152 158218 252847 158454
rect 253083 158218 274916 158454
rect 275152 158218 280847 158454
rect 281083 158218 302916 158454
rect 303152 158218 308847 158454
rect 309083 158218 330916 158454
rect 331152 158218 336847 158454
rect 337083 158218 358916 158454
rect 359152 158218 364847 158454
rect 365083 158218 386916 158454
rect 387152 158218 392847 158454
rect 393083 158218 414916 158454
rect 415152 158218 420847 158454
rect 421083 158218 442916 158454
rect 443152 158218 448847 158454
rect 449083 158218 470916 158454
rect 471152 158218 476847 158454
rect 477083 158218 498916 158454
rect 499152 158218 504847 158454
rect 505083 158218 526916 158454
rect 527152 158218 532847 158454
rect 533083 158218 554916 158454
rect 555152 158218 560847 158454
rect 561083 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 592650 158454
rect -8726 158134 592650 158218
rect -8726 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 22916 158134
rect 23152 157898 28847 158134
rect 29083 157898 50916 158134
rect 51152 157898 56847 158134
rect 57083 157898 78916 158134
rect 79152 157898 84847 158134
rect 85083 157898 106916 158134
rect 107152 157898 112847 158134
rect 113083 157898 134916 158134
rect 135152 157898 140847 158134
rect 141083 157898 162916 158134
rect 163152 157898 168847 158134
rect 169083 157898 190916 158134
rect 191152 157898 196847 158134
rect 197083 157898 218916 158134
rect 219152 157898 224847 158134
rect 225083 157898 246916 158134
rect 247152 157898 252847 158134
rect 253083 157898 274916 158134
rect 275152 157898 280847 158134
rect 281083 157898 302916 158134
rect 303152 157898 308847 158134
rect 309083 157898 330916 158134
rect 331152 157898 336847 158134
rect 337083 157898 358916 158134
rect 359152 157898 364847 158134
rect 365083 157898 386916 158134
rect 387152 157898 392847 158134
rect 393083 157898 414916 158134
rect 415152 157898 420847 158134
rect 421083 157898 442916 158134
rect 443152 157898 448847 158134
rect 449083 157898 470916 158134
rect 471152 157898 476847 158134
rect 477083 157898 498916 158134
rect 499152 157898 504847 158134
rect 505083 157898 526916 158134
rect 527152 157898 532847 158134
rect 533083 157898 554916 158134
rect 555152 157898 560847 158134
rect 561083 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 592650 158134
rect -8726 157866 592650 157898
rect -8726 134829 592650 134861
rect -8726 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 19952 134829
rect 20188 134593 25882 134829
rect 26118 134593 31813 134829
rect 32049 134593 47952 134829
rect 48188 134593 53882 134829
rect 54118 134593 59813 134829
rect 60049 134593 75952 134829
rect 76188 134593 81882 134829
rect 82118 134593 87813 134829
rect 88049 134593 103952 134829
rect 104188 134593 109882 134829
rect 110118 134593 115813 134829
rect 116049 134593 131952 134829
rect 132188 134593 137882 134829
rect 138118 134593 143813 134829
rect 144049 134593 159952 134829
rect 160188 134593 165882 134829
rect 166118 134593 171813 134829
rect 172049 134593 187952 134829
rect 188188 134593 193882 134829
rect 194118 134593 199813 134829
rect 200049 134593 215952 134829
rect 216188 134593 221882 134829
rect 222118 134593 227813 134829
rect 228049 134593 243952 134829
rect 244188 134593 249882 134829
rect 250118 134593 255813 134829
rect 256049 134593 271952 134829
rect 272188 134593 277882 134829
rect 278118 134593 283813 134829
rect 284049 134593 299952 134829
rect 300188 134593 305882 134829
rect 306118 134593 311813 134829
rect 312049 134593 327952 134829
rect 328188 134593 333882 134829
rect 334118 134593 339813 134829
rect 340049 134593 355952 134829
rect 356188 134593 361882 134829
rect 362118 134593 367813 134829
rect 368049 134593 383952 134829
rect 384188 134593 389882 134829
rect 390118 134593 395813 134829
rect 396049 134593 411952 134829
rect 412188 134593 417882 134829
rect 418118 134593 423813 134829
rect 424049 134593 439952 134829
rect 440188 134593 445882 134829
rect 446118 134593 451813 134829
rect 452049 134593 467952 134829
rect 468188 134593 473882 134829
rect 474118 134593 479813 134829
rect 480049 134593 495952 134829
rect 496188 134593 501882 134829
rect 502118 134593 507813 134829
rect 508049 134593 523952 134829
rect 524188 134593 529882 134829
rect 530118 134593 535813 134829
rect 536049 134593 551952 134829
rect 552188 134593 557882 134829
rect 558118 134593 563813 134829
rect 564049 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 592650 134829
rect -8726 134509 592650 134593
rect -8726 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 19952 134509
rect 20188 134273 25882 134509
rect 26118 134273 31813 134509
rect 32049 134273 47952 134509
rect 48188 134273 53882 134509
rect 54118 134273 59813 134509
rect 60049 134273 75952 134509
rect 76188 134273 81882 134509
rect 82118 134273 87813 134509
rect 88049 134273 103952 134509
rect 104188 134273 109882 134509
rect 110118 134273 115813 134509
rect 116049 134273 131952 134509
rect 132188 134273 137882 134509
rect 138118 134273 143813 134509
rect 144049 134273 159952 134509
rect 160188 134273 165882 134509
rect 166118 134273 171813 134509
rect 172049 134273 187952 134509
rect 188188 134273 193882 134509
rect 194118 134273 199813 134509
rect 200049 134273 215952 134509
rect 216188 134273 221882 134509
rect 222118 134273 227813 134509
rect 228049 134273 243952 134509
rect 244188 134273 249882 134509
rect 250118 134273 255813 134509
rect 256049 134273 271952 134509
rect 272188 134273 277882 134509
rect 278118 134273 283813 134509
rect 284049 134273 299952 134509
rect 300188 134273 305882 134509
rect 306118 134273 311813 134509
rect 312049 134273 327952 134509
rect 328188 134273 333882 134509
rect 334118 134273 339813 134509
rect 340049 134273 355952 134509
rect 356188 134273 361882 134509
rect 362118 134273 367813 134509
rect 368049 134273 383952 134509
rect 384188 134273 389882 134509
rect 390118 134273 395813 134509
rect 396049 134273 411952 134509
rect 412188 134273 417882 134509
rect 418118 134273 423813 134509
rect 424049 134273 439952 134509
rect 440188 134273 445882 134509
rect 446118 134273 451813 134509
rect 452049 134273 467952 134509
rect 468188 134273 473882 134509
rect 474118 134273 479813 134509
rect 480049 134273 495952 134509
rect 496188 134273 501882 134509
rect 502118 134273 507813 134509
rect 508049 134273 523952 134509
rect 524188 134273 529882 134509
rect 530118 134273 535813 134509
rect 536049 134273 551952 134509
rect 552188 134273 557882 134509
rect 558118 134273 563813 134509
rect 564049 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 592650 134509
rect -8726 134241 592650 134273
rect -8726 131454 592650 131486
rect -8726 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 22916 131454
rect 23152 131218 28847 131454
rect 29083 131218 50916 131454
rect 51152 131218 56847 131454
rect 57083 131218 78916 131454
rect 79152 131218 84847 131454
rect 85083 131218 106916 131454
rect 107152 131218 112847 131454
rect 113083 131218 134916 131454
rect 135152 131218 140847 131454
rect 141083 131218 162916 131454
rect 163152 131218 168847 131454
rect 169083 131218 190916 131454
rect 191152 131218 196847 131454
rect 197083 131218 218916 131454
rect 219152 131218 224847 131454
rect 225083 131218 246916 131454
rect 247152 131218 252847 131454
rect 253083 131218 274916 131454
rect 275152 131218 280847 131454
rect 281083 131218 302916 131454
rect 303152 131218 308847 131454
rect 309083 131218 330916 131454
rect 331152 131218 336847 131454
rect 337083 131218 358916 131454
rect 359152 131218 364847 131454
rect 365083 131218 386916 131454
rect 387152 131218 392847 131454
rect 393083 131218 414916 131454
rect 415152 131218 420847 131454
rect 421083 131218 442916 131454
rect 443152 131218 448847 131454
rect 449083 131218 470916 131454
rect 471152 131218 476847 131454
rect 477083 131218 498916 131454
rect 499152 131218 504847 131454
rect 505083 131218 526916 131454
rect 527152 131218 532847 131454
rect 533083 131218 554916 131454
rect 555152 131218 560847 131454
rect 561083 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 592650 131454
rect -8726 131134 592650 131218
rect -8726 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 22916 131134
rect 23152 130898 28847 131134
rect 29083 130898 50916 131134
rect 51152 130898 56847 131134
rect 57083 130898 78916 131134
rect 79152 130898 84847 131134
rect 85083 130898 106916 131134
rect 107152 130898 112847 131134
rect 113083 130898 134916 131134
rect 135152 130898 140847 131134
rect 141083 130898 162916 131134
rect 163152 130898 168847 131134
rect 169083 130898 190916 131134
rect 191152 130898 196847 131134
rect 197083 130898 218916 131134
rect 219152 130898 224847 131134
rect 225083 130898 246916 131134
rect 247152 130898 252847 131134
rect 253083 130898 274916 131134
rect 275152 130898 280847 131134
rect 281083 130898 302916 131134
rect 303152 130898 308847 131134
rect 309083 130898 330916 131134
rect 331152 130898 336847 131134
rect 337083 130898 358916 131134
rect 359152 130898 364847 131134
rect 365083 130898 386916 131134
rect 387152 130898 392847 131134
rect 393083 130898 414916 131134
rect 415152 130898 420847 131134
rect 421083 130898 442916 131134
rect 443152 130898 448847 131134
rect 449083 130898 470916 131134
rect 471152 130898 476847 131134
rect 477083 130898 498916 131134
rect 499152 130898 504847 131134
rect 505083 130898 526916 131134
rect 527152 130898 532847 131134
rect 533083 130898 554916 131134
rect 555152 130898 560847 131134
rect 561083 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 592650 131134
rect -8726 130866 592650 130898
rect -8726 107829 592650 107861
rect -8726 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 19952 107829
rect 20188 107593 25882 107829
rect 26118 107593 31813 107829
rect 32049 107593 47952 107829
rect 48188 107593 53882 107829
rect 54118 107593 59813 107829
rect 60049 107593 75952 107829
rect 76188 107593 81882 107829
rect 82118 107593 87813 107829
rect 88049 107593 103952 107829
rect 104188 107593 109882 107829
rect 110118 107593 115813 107829
rect 116049 107593 131952 107829
rect 132188 107593 137882 107829
rect 138118 107593 143813 107829
rect 144049 107593 159952 107829
rect 160188 107593 165882 107829
rect 166118 107593 171813 107829
rect 172049 107593 187952 107829
rect 188188 107593 193882 107829
rect 194118 107593 199813 107829
rect 200049 107593 215952 107829
rect 216188 107593 221882 107829
rect 222118 107593 227813 107829
rect 228049 107593 243952 107829
rect 244188 107593 249882 107829
rect 250118 107593 255813 107829
rect 256049 107593 271952 107829
rect 272188 107593 277882 107829
rect 278118 107593 283813 107829
rect 284049 107593 299952 107829
rect 300188 107593 305882 107829
rect 306118 107593 311813 107829
rect 312049 107593 327952 107829
rect 328188 107593 333882 107829
rect 334118 107593 339813 107829
rect 340049 107593 355952 107829
rect 356188 107593 361882 107829
rect 362118 107593 367813 107829
rect 368049 107593 383952 107829
rect 384188 107593 389882 107829
rect 390118 107593 395813 107829
rect 396049 107593 411952 107829
rect 412188 107593 417882 107829
rect 418118 107593 423813 107829
rect 424049 107593 439952 107829
rect 440188 107593 445882 107829
rect 446118 107593 451813 107829
rect 452049 107593 467952 107829
rect 468188 107593 473882 107829
rect 474118 107593 479813 107829
rect 480049 107593 495952 107829
rect 496188 107593 501882 107829
rect 502118 107593 507813 107829
rect 508049 107593 523952 107829
rect 524188 107593 529882 107829
rect 530118 107593 535813 107829
rect 536049 107593 551952 107829
rect 552188 107593 557882 107829
rect 558118 107593 563813 107829
rect 564049 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 592650 107829
rect -8726 107509 592650 107593
rect -8726 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 19952 107509
rect 20188 107273 25882 107509
rect 26118 107273 31813 107509
rect 32049 107273 47952 107509
rect 48188 107273 53882 107509
rect 54118 107273 59813 107509
rect 60049 107273 75952 107509
rect 76188 107273 81882 107509
rect 82118 107273 87813 107509
rect 88049 107273 103952 107509
rect 104188 107273 109882 107509
rect 110118 107273 115813 107509
rect 116049 107273 131952 107509
rect 132188 107273 137882 107509
rect 138118 107273 143813 107509
rect 144049 107273 159952 107509
rect 160188 107273 165882 107509
rect 166118 107273 171813 107509
rect 172049 107273 187952 107509
rect 188188 107273 193882 107509
rect 194118 107273 199813 107509
rect 200049 107273 215952 107509
rect 216188 107273 221882 107509
rect 222118 107273 227813 107509
rect 228049 107273 243952 107509
rect 244188 107273 249882 107509
rect 250118 107273 255813 107509
rect 256049 107273 271952 107509
rect 272188 107273 277882 107509
rect 278118 107273 283813 107509
rect 284049 107273 299952 107509
rect 300188 107273 305882 107509
rect 306118 107273 311813 107509
rect 312049 107273 327952 107509
rect 328188 107273 333882 107509
rect 334118 107273 339813 107509
rect 340049 107273 355952 107509
rect 356188 107273 361882 107509
rect 362118 107273 367813 107509
rect 368049 107273 383952 107509
rect 384188 107273 389882 107509
rect 390118 107273 395813 107509
rect 396049 107273 411952 107509
rect 412188 107273 417882 107509
rect 418118 107273 423813 107509
rect 424049 107273 439952 107509
rect 440188 107273 445882 107509
rect 446118 107273 451813 107509
rect 452049 107273 467952 107509
rect 468188 107273 473882 107509
rect 474118 107273 479813 107509
rect 480049 107273 495952 107509
rect 496188 107273 501882 107509
rect 502118 107273 507813 107509
rect 508049 107273 523952 107509
rect 524188 107273 529882 107509
rect 530118 107273 535813 107509
rect 536049 107273 551952 107509
rect 552188 107273 557882 107509
rect 558118 107273 563813 107509
rect 564049 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 592650 107509
rect -8726 107241 592650 107273
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 22916 104454
rect 23152 104218 28847 104454
rect 29083 104218 50916 104454
rect 51152 104218 56847 104454
rect 57083 104218 78916 104454
rect 79152 104218 84847 104454
rect 85083 104218 106916 104454
rect 107152 104218 112847 104454
rect 113083 104218 134916 104454
rect 135152 104218 140847 104454
rect 141083 104218 162916 104454
rect 163152 104218 168847 104454
rect 169083 104218 190916 104454
rect 191152 104218 196847 104454
rect 197083 104218 218916 104454
rect 219152 104218 224847 104454
rect 225083 104218 246916 104454
rect 247152 104218 252847 104454
rect 253083 104218 274916 104454
rect 275152 104218 280847 104454
rect 281083 104218 302916 104454
rect 303152 104218 308847 104454
rect 309083 104218 330916 104454
rect 331152 104218 336847 104454
rect 337083 104218 358916 104454
rect 359152 104218 364847 104454
rect 365083 104218 386916 104454
rect 387152 104218 392847 104454
rect 393083 104218 414916 104454
rect 415152 104218 420847 104454
rect 421083 104218 442916 104454
rect 443152 104218 448847 104454
rect 449083 104218 470916 104454
rect 471152 104218 476847 104454
rect 477083 104218 498916 104454
rect 499152 104218 504847 104454
rect 505083 104218 526916 104454
rect 527152 104218 532847 104454
rect 533083 104218 554916 104454
rect 555152 104218 560847 104454
rect 561083 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 22916 104134
rect 23152 103898 28847 104134
rect 29083 103898 50916 104134
rect 51152 103898 56847 104134
rect 57083 103898 78916 104134
rect 79152 103898 84847 104134
rect 85083 103898 106916 104134
rect 107152 103898 112847 104134
rect 113083 103898 134916 104134
rect 135152 103898 140847 104134
rect 141083 103898 162916 104134
rect 163152 103898 168847 104134
rect 169083 103898 190916 104134
rect 191152 103898 196847 104134
rect 197083 103898 218916 104134
rect 219152 103898 224847 104134
rect 225083 103898 246916 104134
rect 247152 103898 252847 104134
rect 253083 103898 274916 104134
rect 275152 103898 280847 104134
rect 281083 103898 302916 104134
rect 303152 103898 308847 104134
rect 309083 103898 330916 104134
rect 331152 103898 336847 104134
rect 337083 103898 358916 104134
rect 359152 103898 364847 104134
rect 365083 103898 386916 104134
rect 387152 103898 392847 104134
rect 393083 103898 414916 104134
rect 415152 103898 420847 104134
rect 421083 103898 442916 104134
rect 443152 103898 448847 104134
rect 449083 103898 470916 104134
rect 471152 103898 476847 104134
rect 477083 103898 498916 104134
rect 499152 103898 504847 104134
rect 505083 103898 526916 104134
rect 527152 103898 532847 104134
rect 533083 103898 554916 104134
rect 555152 103898 560847 104134
rect 561083 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 80829 592650 80861
rect -8726 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 19952 80829
rect 20188 80593 25882 80829
rect 26118 80593 31813 80829
rect 32049 80593 47952 80829
rect 48188 80593 53882 80829
rect 54118 80593 59813 80829
rect 60049 80593 75952 80829
rect 76188 80593 81882 80829
rect 82118 80593 87813 80829
rect 88049 80593 103952 80829
rect 104188 80593 109882 80829
rect 110118 80593 115813 80829
rect 116049 80593 131952 80829
rect 132188 80593 137882 80829
rect 138118 80593 143813 80829
rect 144049 80593 159952 80829
rect 160188 80593 165882 80829
rect 166118 80593 171813 80829
rect 172049 80593 187952 80829
rect 188188 80593 193882 80829
rect 194118 80593 199813 80829
rect 200049 80593 215952 80829
rect 216188 80593 221882 80829
rect 222118 80593 227813 80829
rect 228049 80593 243952 80829
rect 244188 80593 249882 80829
rect 250118 80593 255813 80829
rect 256049 80593 271952 80829
rect 272188 80593 277882 80829
rect 278118 80593 283813 80829
rect 284049 80593 299952 80829
rect 300188 80593 305882 80829
rect 306118 80593 311813 80829
rect 312049 80593 327952 80829
rect 328188 80593 333882 80829
rect 334118 80593 339813 80829
rect 340049 80593 355952 80829
rect 356188 80593 361882 80829
rect 362118 80593 367813 80829
rect 368049 80593 383952 80829
rect 384188 80593 389882 80829
rect 390118 80593 395813 80829
rect 396049 80593 411952 80829
rect 412188 80593 417882 80829
rect 418118 80593 423813 80829
rect 424049 80593 439952 80829
rect 440188 80593 445882 80829
rect 446118 80593 451813 80829
rect 452049 80593 467952 80829
rect 468188 80593 473882 80829
rect 474118 80593 479813 80829
rect 480049 80593 495952 80829
rect 496188 80593 501882 80829
rect 502118 80593 507813 80829
rect 508049 80593 523952 80829
rect 524188 80593 529882 80829
rect 530118 80593 535813 80829
rect 536049 80593 551952 80829
rect 552188 80593 557882 80829
rect 558118 80593 563813 80829
rect 564049 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 592650 80829
rect -8726 80509 592650 80593
rect -8726 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 19952 80509
rect 20188 80273 25882 80509
rect 26118 80273 31813 80509
rect 32049 80273 47952 80509
rect 48188 80273 53882 80509
rect 54118 80273 59813 80509
rect 60049 80273 75952 80509
rect 76188 80273 81882 80509
rect 82118 80273 87813 80509
rect 88049 80273 103952 80509
rect 104188 80273 109882 80509
rect 110118 80273 115813 80509
rect 116049 80273 131952 80509
rect 132188 80273 137882 80509
rect 138118 80273 143813 80509
rect 144049 80273 159952 80509
rect 160188 80273 165882 80509
rect 166118 80273 171813 80509
rect 172049 80273 187952 80509
rect 188188 80273 193882 80509
rect 194118 80273 199813 80509
rect 200049 80273 215952 80509
rect 216188 80273 221882 80509
rect 222118 80273 227813 80509
rect 228049 80273 243952 80509
rect 244188 80273 249882 80509
rect 250118 80273 255813 80509
rect 256049 80273 271952 80509
rect 272188 80273 277882 80509
rect 278118 80273 283813 80509
rect 284049 80273 299952 80509
rect 300188 80273 305882 80509
rect 306118 80273 311813 80509
rect 312049 80273 327952 80509
rect 328188 80273 333882 80509
rect 334118 80273 339813 80509
rect 340049 80273 355952 80509
rect 356188 80273 361882 80509
rect 362118 80273 367813 80509
rect 368049 80273 383952 80509
rect 384188 80273 389882 80509
rect 390118 80273 395813 80509
rect 396049 80273 411952 80509
rect 412188 80273 417882 80509
rect 418118 80273 423813 80509
rect 424049 80273 439952 80509
rect 440188 80273 445882 80509
rect 446118 80273 451813 80509
rect 452049 80273 467952 80509
rect 468188 80273 473882 80509
rect 474118 80273 479813 80509
rect 480049 80273 495952 80509
rect 496188 80273 501882 80509
rect 502118 80273 507813 80509
rect 508049 80273 523952 80509
rect 524188 80273 529882 80509
rect 530118 80273 535813 80509
rect 536049 80273 551952 80509
rect 552188 80273 557882 80509
rect 558118 80273 563813 80509
rect 564049 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 592650 80509
rect -8726 80241 592650 80273
rect -8726 77454 592650 77486
rect -8726 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 22916 77454
rect 23152 77218 28847 77454
rect 29083 77218 50916 77454
rect 51152 77218 56847 77454
rect 57083 77218 78916 77454
rect 79152 77218 84847 77454
rect 85083 77218 106916 77454
rect 107152 77218 112847 77454
rect 113083 77218 134916 77454
rect 135152 77218 140847 77454
rect 141083 77218 162916 77454
rect 163152 77218 168847 77454
rect 169083 77218 190916 77454
rect 191152 77218 196847 77454
rect 197083 77218 218916 77454
rect 219152 77218 224847 77454
rect 225083 77218 246916 77454
rect 247152 77218 252847 77454
rect 253083 77218 274916 77454
rect 275152 77218 280847 77454
rect 281083 77218 302916 77454
rect 303152 77218 308847 77454
rect 309083 77218 330916 77454
rect 331152 77218 336847 77454
rect 337083 77218 358916 77454
rect 359152 77218 364847 77454
rect 365083 77218 386916 77454
rect 387152 77218 392847 77454
rect 393083 77218 414916 77454
rect 415152 77218 420847 77454
rect 421083 77218 442916 77454
rect 443152 77218 448847 77454
rect 449083 77218 470916 77454
rect 471152 77218 476847 77454
rect 477083 77218 498916 77454
rect 499152 77218 504847 77454
rect 505083 77218 526916 77454
rect 527152 77218 532847 77454
rect 533083 77218 554916 77454
rect 555152 77218 560847 77454
rect 561083 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 592650 77454
rect -8726 77134 592650 77218
rect -8726 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 22916 77134
rect 23152 76898 28847 77134
rect 29083 76898 50916 77134
rect 51152 76898 56847 77134
rect 57083 76898 78916 77134
rect 79152 76898 84847 77134
rect 85083 76898 106916 77134
rect 107152 76898 112847 77134
rect 113083 76898 134916 77134
rect 135152 76898 140847 77134
rect 141083 76898 162916 77134
rect 163152 76898 168847 77134
rect 169083 76898 190916 77134
rect 191152 76898 196847 77134
rect 197083 76898 218916 77134
rect 219152 76898 224847 77134
rect 225083 76898 246916 77134
rect 247152 76898 252847 77134
rect 253083 76898 274916 77134
rect 275152 76898 280847 77134
rect 281083 76898 302916 77134
rect 303152 76898 308847 77134
rect 309083 76898 330916 77134
rect 331152 76898 336847 77134
rect 337083 76898 358916 77134
rect 359152 76898 364847 77134
rect 365083 76898 386916 77134
rect 387152 76898 392847 77134
rect 393083 76898 414916 77134
rect 415152 76898 420847 77134
rect 421083 76898 442916 77134
rect 443152 76898 448847 77134
rect 449083 76898 470916 77134
rect 471152 76898 476847 77134
rect 477083 76898 498916 77134
rect 499152 76898 504847 77134
rect 505083 76898 526916 77134
rect 527152 76898 532847 77134
rect 533083 76898 554916 77134
rect 555152 76898 560847 77134
rect 561083 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 592650 77134
rect -8726 76866 592650 76898
rect -8726 53829 592650 53861
rect -8726 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 19952 53829
rect 20188 53593 25882 53829
rect 26118 53593 31813 53829
rect 32049 53593 47952 53829
rect 48188 53593 53882 53829
rect 54118 53593 59813 53829
rect 60049 53593 75952 53829
rect 76188 53593 81882 53829
rect 82118 53593 87813 53829
rect 88049 53593 103952 53829
rect 104188 53593 109882 53829
rect 110118 53593 115813 53829
rect 116049 53593 131952 53829
rect 132188 53593 137882 53829
rect 138118 53593 143813 53829
rect 144049 53593 159952 53829
rect 160188 53593 165882 53829
rect 166118 53593 171813 53829
rect 172049 53593 187952 53829
rect 188188 53593 193882 53829
rect 194118 53593 199813 53829
rect 200049 53593 215952 53829
rect 216188 53593 221882 53829
rect 222118 53593 227813 53829
rect 228049 53593 243952 53829
rect 244188 53593 249882 53829
rect 250118 53593 255813 53829
rect 256049 53593 271952 53829
rect 272188 53593 277882 53829
rect 278118 53593 283813 53829
rect 284049 53593 299952 53829
rect 300188 53593 305882 53829
rect 306118 53593 311813 53829
rect 312049 53593 327952 53829
rect 328188 53593 333882 53829
rect 334118 53593 339813 53829
rect 340049 53593 355952 53829
rect 356188 53593 361882 53829
rect 362118 53593 367813 53829
rect 368049 53593 383952 53829
rect 384188 53593 389882 53829
rect 390118 53593 395813 53829
rect 396049 53593 411952 53829
rect 412188 53593 417882 53829
rect 418118 53593 423813 53829
rect 424049 53593 439952 53829
rect 440188 53593 445882 53829
rect 446118 53593 451813 53829
rect 452049 53593 467952 53829
rect 468188 53593 473882 53829
rect 474118 53593 479813 53829
rect 480049 53593 495952 53829
rect 496188 53593 501882 53829
rect 502118 53593 507813 53829
rect 508049 53593 523952 53829
rect 524188 53593 529882 53829
rect 530118 53593 535813 53829
rect 536049 53593 551952 53829
rect 552188 53593 557882 53829
rect 558118 53593 563813 53829
rect 564049 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 592650 53829
rect -8726 53509 592650 53593
rect -8726 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 19952 53509
rect 20188 53273 25882 53509
rect 26118 53273 31813 53509
rect 32049 53273 47952 53509
rect 48188 53273 53882 53509
rect 54118 53273 59813 53509
rect 60049 53273 75952 53509
rect 76188 53273 81882 53509
rect 82118 53273 87813 53509
rect 88049 53273 103952 53509
rect 104188 53273 109882 53509
rect 110118 53273 115813 53509
rect 116049 53273 131952 53509
rect 132188 53273 137882 53509
rect 138118 53273 143813 53509
rect 144049 53273 159952 53509
rect 160188 53273 165882 53509
rect 166118 53273 171813 53509
rect 172049 53273 187952 53509
rect 188188 53273 193882 53509
rect 194118 53273 199813 53509
rect 200049 53273 215952 53509
rect 216188 53273 221882 53509
rect 222118 53273 227813 53509
rect 228049 53273 243952 53509
rect 244188 53273 249882 53509
rect 250118 53273 255813 53509
rect 256049 53273 271952 53509
rect 272188 53273 277882 53509
rect 278118 53273 283813 53509
rect 284049 53273 299952 53509
rect 300188 53273 305882 53509
rect 306118 53273 311813 53509
rect 312049 53273 327952 53509
rect 328188 53273 333882 53509
rect 334118 53273 339813 53509
rect 340049 53273 355952 53509
rect 356188 53273 361882 53509
rect 362118 53273 367813 53509
rect 368049 53273 383952 53509
rect 384188 53273 389882 53509
rect 390118 53273 395813 53509
rect 396049 53273 411952 53509
rect 412188 53273 417882 53509
rect 418118 53273 423813 53509
rect 424049 53273 439952 53509
rect 440188 53273 445882 53509
rect 446118 53273 451813 53509
rect 452049 53273 467952 53509
rect 468188 53273 473882 53509
rect 474118 53273 479813 53509
rect 480049 53273 495952 53509
rect 496188 53273 501882 53509
rect 502118 53273 507813 53509
rect 508049 53273 523952 53509
rect 524188 53273 529882 53509
rect 530118 53273 535813 53509
rect 536049 53273 551952 53509
rect 552188 53273 557882 53509
rect 558118 53273 563813 53509
rect 564049 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 592650 53509
rect -8726 53241 592650 53273
rect -8726 50454 592650 50486
rect -8726 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 22916 50454
rect 23152 50218 28847 50454
rect 29083 50218 50916 50454
rect 51152 50218 56847 50454
rect 57083 50218 78916 50454
rect 79152 50218 84847 50454
rect 85083 50218 106916 50454
rect 107152 50218 112847 50454
rect 113083 50218 134916 50454
rect 135152 50218 140847 50454
rect 141083 50218 162916 50454
rect 163152 50218 168847 50454
rect 169083 50218 190916 50454
rect 191152 50218 196847 50454
rect 197083 50218 218916 50454
rect 219152 50218 224847 50454
rect 225083 50218 246916 50454
rect 247152 50218 252847 50454
rect 253083 50218 274916 50454
rect 275152 50218 280847 50454
rect 281083 50218 302916 50454
rect 303152 50218 308847 50454
rect 309083 50218 330916 50454
rect 331152 50218 336847 50454
rect 337083 50218 358916 50454
rect 359152 50218 364847 50454
rect 365083 50218 386916 50454
rect 387152 50218 392847 50454
rect 393083 50218 414916 50454
rect 415152 50218 420847 50454
rect 421083 50218 442916 50454
rect 443152 50218 448847 50454
rect 449083 50218 470916 50454
rect 471152 50218 476847 50454
rect 477083 50218 498916 50454
rect 499152 50218 504847 50454
rect 505083 50218 526916 50454
rect 527152 50218 532847 50454
rect 533083 50218 554916 50454
rect 555152 50218 560847 50454
rect 561083 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 592650 50454
rect -8726 50134 592650 50218
rect -8726 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 22916 50134
rect 23152 49898 28847 50134
rect 29083 49898 50916 50134
rect 51152 49898 56847 50134
rect 57083 49898 78916 50134
rect 79152 49898 84847 50134
rect 85083 49898 106916 50134
rect 107152 49898 112847 50134
rect 113083 49898 134916 50134
rect 135152 49898 140847 50134
rect 141083 49898 162916 50134
rect 163152 49898 168847 50134
rect 169083 49898 190916 50134
rect 191152 49898 196847 50134
rect 197083 49898 218916 50134
rect 219152 49898 224847 50134
rect 225083 49898 246916 50134
rect 247152 49898 252847 50134
rect 253083 49898 274916 50134
rect 275152 49898 280847 50134
rect 281083 49898 302916 50134
rect 303152 49898 308847 50134
rect 309083 49898 330916 50134
rect 331152 49898 336847 50134
rect 337083 49898 358916 50134
rect 359152 49898 364847 50134
rect 365083 49898 386916 50134
rect 387152 49898 392847 50134
rect 393083 49898 414916 50134
rect 415152 49898 420847 50134
rect 421083 49898 442916 50134
rect 443152 49898 448847 50134
rect 449083 49898 470916 50134
rect 471152 49898 476847 50134
rect 477083 49898 498916 50134
rect 499152 49898 504847 50134
rect 505083 49898 526916 50134
rect 527152 49898 532847 50134
rect 533083 49898 554916 50134
rect 555152 49898 560847 50134
rect 561083 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 592650 50134
rect -8726 49866 592650 49898
rect -8726 26829 592650 26861
rect -8726 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 24284 26829
rect 24520 26593 38882 26829
rect 39118 26593 53479 26829
rect 53715 26593 75952 26829
rect 76188 26593 81882 26829
rect 82118 26593 87813 26829
rect 88049 26593 103952 26829
rect 104188 26593 109882 26829
rect 110118 26593 115813 26829
rect 116049 26593 131952 26829
rect 132188 26593 137882 26829
rect 138118 26593 143813 26829
rect 144049 26593 159952 26829
rect 160188 26593 165882 26829
rect 166118 26593 171813 26829
rect 172049 26593 187952 26829
rect 188188 26593 193882 26829
rect 194118 26593 199813 26829
rect 200049 26593 215952 26829
rect 216188 26593 221882 26829
rect 222118 26593 227813 26829
rect 228049 26593 243952 26829
rect 244188 26593 249882 26829
rect 250118 26593 255813 26829
rect 256049 26593 271952 26829
rect 272188 26593 277882 26829
rect 278118 26593 283813 26829
rect 284049 26593 299952 26829
rect 300188 26593 305882 26829
rect 306118 26593 311813 26829
rect 312049 26593 327952 26829
rect 328188 26593 333882 26829
rect 334118 26593 339813 26829
rect 340049 26593 355952 26829
rect 356188 26593 361882 26829
rect 362118 26593 367813 26829
rect 368049 26593 383952 26829
rect 384188 26593 389882 26829
rect 390118 26593 395813 26829
rect 396049 26593 411952 26829
rect 412188 26593 417882 26829
rect 418118 26593 423813 26829
rect 424049 26593 439952 26829
rect 440188 26593 445882 26829
rect 446118 26593 451813 26829
rect 452049 26593 467952 26829
rect 468188 26593 473882 26829
rect 474118 26593 479813 26829
rect 480049 26593 495952 26829
rect 496188 26593 501882 26829
rect 502118 26593 507813 26829
rect 508049 26593 523952 26829
rect 524188 26593 529882 26829
rect 530118 26593 535813 26829
rect 536049 26593 551952 26829
rect 552188 26593 557882 26829
rect 558118 26593 563813 26829
rect 564049 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 592650 26829
rect -8726 26509 592650 26593
rect -8726 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 24284 26509
rect 24520 26273 38882 26509
rect 39118 26273 53479 26509
rect 53715 26273 75952 26509
rect 76188 26273 81882 26509
rect 82118 26273 87813 26509
rect 88049 26273 103952 26509
rect 104188 26273 109882 26509
rect 110118 26273 115813 26509
rect 116049 26273 131952 26509
rect 132188 26273 137882 26509
rect 138118 26273 143813 26509
rect 144049 26273 159952 26509
rect 160188 26273 165882 26509
rect 166118 26273 171813 26509
rect 172049 26273 187952 26509
rect 188188 26273 193882 26509
rect 194118 26273 199813 26509
rect 200049 26273 215952 26509
rect 216188 26273 221882 26509
rect 222118 26273 227813 26509
rect 228049 26273 243952 26509
rect 244188 26273 249882 26509
rect 250118 26273 255813 26509
rect 256049 26273 271952 26509
rect 272188 26273 277882 26509
rect 278118 26273 283813 26509
rect 284049 26273 299952 26509
rect 300188 26273 305882 26509
rect 306118 26273 311813 26509
rect 312049 26273 327952 26509
rect 328188 26273 333882 26509
rect 334118 26273 339813 26509
rect 340049 26273 355952 26509
rect 356188 26273 361882 26509
rect 362118 26273 367813 26509
rect 368049 26273 383952 26509
rect 384188 26273 389882 26509
rect 390118 26273 395813 26509
rect 396049 26273 411952 26509
rect 412188 26273 417882 26509
rect 418118 26273 423813 26509
rect 424049 26273 439952 26509
rect 440188 26273 445882 26509
rect 446118 26273 451813 26509
rect 452049 26273 467952 26509
rect 468188 26273 473882 26509
rect 474118 26273 479813 26509
rect 480049 26273 495952 26509
rect 496188 26273 501882 26509
rect 502118 26273 507813 26509
rect 508049 26273 523952 26509
rect 524188 26273 529882 26509
rect 530118 26273 535813 26509
rect 536049 26273 551952 26509
rect 552188 26273 557882 26509
rect 558118 26273 563813 26509
rect 564049 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 592650 26509
rect -8726 26241 592650 26273
rect -8726 23454 592650 23486
rect -8726 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 31584 23454
rect 31820 23218 46181 23454
rect 46417 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 78916 23454
rect 79152 23218 84847 23454
rect 85083 23218 106916 23454
rect 107152 23218 112847 23454
rect 113083 23218 134916 23454
rect 135152 23218 140847 23454
rect 141083 23218 162916 23454
rect 163152 23218 168847 23454
rect 169083 23218 190916 23454
rect 191152 23218 196847 23454
rect 197083 23218 218916 23454
rect 219152 23218 224847 23454
rect 225083 23218 246916 23454
rect 247152 23218 252847 23454
rect 253083 23218 274916 23454
rect 275152 23218 280847 23454
rect 281083 23218 302916 23454
rect 303152 23218 308847 23454
rect 309083 23218 330916 23454
rect 331152 23218 336847 23454
rect 337083 23218 358916 23454
rect 359152 23218 364847 23454
rect 365083 23218 386916 23454
rect 387152 23218 392847 23454
rect 393083 23218 414916 23454
rect 415152 23218 420847 23454
rect 421083 23218 442916 23454
rect 443152 23218 448847 23454
rect 449083 23218 470916 23454
rect 471152 23218 476847 23454
rect 477083 23218 498916 23454
rect 499152 23218 504847 23454
rect 505083 23218 526916 23454
rect 527152 23218 532847 23454
rect 533083 23218 554916 23454
rect 555152 23218 560847 23454
rect 561083 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 592650 23454
rect -8726 23134 592650 23218
rect -8726 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 31584 23134
rect 31820 22898 46181 23134
rect 46417 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 78916 23134
rect 79152 22898 84847 23134
rect 85083 22898 106916 23134
rect 107152 22898 112847 23134
rect 113083 22898 134916 23134
rect 135152 22898 140847 23134
rect 141083 22898 162916 23134
rect 163152 22898 168847 23134
rect 169083 22898 190916 23134
rect 191152 22898 196847 23134
rect 197083 22898 218916 23134
rect 219152 22898 224847 23134
rect 225083 22898 246916 23134
rect 247152 22898 252847 23134
rect 253083 22898 274916 23134
rect 275152 22898 280847 23134
rect 281083 22898 302916 23134
rect 303152 22898 308847 23134
rect 309083 22898 330916 23134
rect 331152 22898 336847 23134
rect 337083 22898 358916 23134
rect 359152 22898 364847 23134
rect 365083 22898 386916 23134
rect 387152 22898 392847 23134
rect 393083 22898 414916 23134
rect 415152 22898 420847 23134
rect 421083 22898 442916 23134
rect 443152 22898 448847 23134
rect 449083 22898 470916 23134
rect 471152 22898 476847 23134
rect 477083 22898 498916 23134
rect 499152 22898 504847 23134
rect 505083 22898 526916 23134
rect 527152 22898 532847 23134
rect 533083 22898 554916 23134
rect 555152 22898 560847 23134
rect 561083 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 592650 23134
rect -8726 22866 592650 22898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use scan_controller  scan_controller
timestamp 0
transform 1 0 16000 0 1 16000
box -10 -52 46000 20000
use scan_wrapper_334445762078310996  scan_wrapper_334445762078310996_1
timestamp 0
transform 1 0 100000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_335404063203000914  scan_wrapper_335404063203000914_2
timestamp 0
transform 1 0 128000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339439899388150354  scan_wrapper_339439899388150354_3
timestamp 0
transform 1 0 156000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_0
timestamp 0
transform 1 0 72000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_13
timestamp 0
transform 1 0 436000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_14
timestamp 0
transform 1 0 464000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_15
timestamp 0
transform 1 0 492000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_16
timestamp 0
transform 1 0 520000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_17
timestamp 0
transform 1 0 548000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_18
timestamp 0
transform 1 0 16000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_19
timestamp 0
transform 1 0 44000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_20
timestamp 0
transform 1 0 72000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_21
timestamp 0
transform 1 0 100000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_22
timestamp 0
transform 1 0 128000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_23
timestamp 0
transform 1 0 156000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_24
timestamp 0
transform 1 0 184000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_25
timestamp 0
transform 1 0 212000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_26
timestamp 0
transform 1 0 240000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_27
timestamp 0
transform 1 0 268000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_28
timestamp 0
transform 1 0 296000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_29
timestamp 0
transform 1 0 324000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_30
timestamp 0
transform 1 0 352000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_31
timestamp 0
transform 1 0 380000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_32
timestamp 0
transform 1 0 408000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_33
timestamp 0
transform 1 0 436000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_34
timestamp 0
transform 1 0 464000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_35
timestamp 0
transform 1 0 492000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_36
timestamp 0
transform 1 0 520000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_37
timestamp 0
transform 1 0 548000 0 1 43000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_38
timestamp 0
transform 1 0 16000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_39
timestamp 0
transform 1 0 44000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_40
timestamp 0
transform 1 0 72000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_41
timestamp 0
transform 1 0 100000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_42
timestamp 0
transform 1 0 128000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_43
timestamp 0
transform 1 0 156000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_44
timestamp 0
transform 1 0 184000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_45
timestamp 0
transform 1 0 212000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_46
timestamp 0
transform 1 0 240000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_47
timestamp 0
transform 1 0 268000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_48
timestamp 0
transform 1 0 296000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_49
timestamp 0
transform 1 0 324000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_50
timestamp 0
transform 1 0 352000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_51
timestamp 0
transform 1 0 380000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_52
timestamp 0
transform 1 0 408000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_53
timestamp 0
transform 1 0 436000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_54
timestamp 0
transform 1 0 464000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_55
timestamp 0
transform 1 0 492000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_56
timestamp 0
transform 1 0 520000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_57
timestamp 0
transform 1 0 548000 0 1 70000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_58
timestamp 0
transform 1 0 16000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_59
timestamp 0
transform 1 0 44000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_60
timestamp 0
transform 1 0 72000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_61
timestamp 0
transform 1 0 100000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_62
timestamp 0
transform 1 0 128000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_63
timestamp 0
transform 1 0 156000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_64
timestamp 0
transform 1 0 184000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_65
timestamp 0
transform 1 0 212000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_66
timestamp 0
transform 1 0 240000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_67
timestamp 0
transform 1 0 268000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_68
timestamp 0
transform 1 0 296000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_69
timestamp 0
transform 1 0 324000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_70
timestamp 0
transform 1 0 352000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_71
timestamp 0
transform 1 0 380000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_72
timestamp 0
transform 1 0 408000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_73
timestamp 0
transform 1 0 436000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_74
timestamp 0
transform 1 0 464000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_75
timestamp 0
transform 1 0 492000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_76
timestamp 0
transform 1 0 520000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_77
timestamp 0
transform 1 0 548000 0 1 97000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_78
timestamp 0
transform 1 0 16000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_79
timestamp 0
transform 1 0 44000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_80
timestamp 0
transform 1 0 72000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_81
timestamp 0
transform 1 0 100000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_82
timestamp 0
transform 1 0 128000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_83
timestamp 0
transform 1 0 156000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_84
timestamp 0
transform 1 0 184000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_85
timestamp 0
transform 1 0 212000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_86
timestamp 0
transform 1 0 240000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_87
timestamp 0
transform 1 0 268000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_88
timestamp 0
transform 1 0 296000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_89
timestamp 0
transform 1 0 324000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_90
timestamp 0
transform 1 0 352000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_91
timestamp 0
transform 1 0 380000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_92
timestamp 0
transform 1 0 408000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_93
timestamp 0
transform 1 0 436000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_94
timestamp 0
transform 1 0 464000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_95
timestamp 0
transform 1 0 492000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_96
timestamp 0
transform 1 0 520000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_97
timestamp 0
transform 1 0 548000 0 1 124000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_98
timestamp 0
transform 1 0 16000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_99
timestamp 0
transform 1 0 44000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_100
timestamp 0
transform 1 0 72000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_101
timestamp 0
transform 1 0 100000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_102
timestamp 0
transform 1 0 128000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_103
timestamp 0
transform 1 0 156000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_104
timestamp 0
transform 1 0 184000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_105
timestamp 0
transform 1 0 212000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_106
timestamp 0
transform 1 0 240000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_107
timestamp 0
transform 1 0 268000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_108
timestamp 0
transform 1 0 296000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_109
timestamp 0
transform 1 0 324000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_110
timestamp 0
transform 1 0 352000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_111
timestamp 0
transform 1 0 380000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_112
timestamp 0
transform 1 0 408000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_113
timestamp 0
transform 1 0 436000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_114
timestamp 0
transform 1 0 464000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_115
timestamp 0
transform 1 0 492000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_116
timestamp 0
transform 1 0 520000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_117
timestamp 0
transform 1 0 548000 0 1 151000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_118
timestamp 0
transform 1 0 16000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_119
timestamp 0
transform 1 0 44000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_120
timestamp 0
transform 1 0 72000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_121
timestamp 0
transform 1 0 100000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_122
timestamp 0
transform 1 0 128000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_123
timestamp 0
transform 1 0 156000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_124
timestamp 0
transform 1 0 184000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_125
timestamp 0
transform 1 0 212000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_126
timestamp 0
transform 1 0 240000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_127
timestamp 0
transform 1 0 268000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_128
timestamp 0
transform 1 0 296000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_129
timestamp 0
transform 1 0 324000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_130
timestamp 0
transform 1 0 352000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_131
timestamp 0
transform 1 0 380000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_132
timestamp 0
transform 1 0 408000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_133
timestamp 0
transform 1 0 436000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_134
timestamp 0
transform 1 0 464000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_135
timestamp 0
transform 1 0 492000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_136
timestamp 0
transform 1 0 520000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_137
timestamp 0
transform 1 0 548000 0 1 178000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_138
timestamp 0
transform 1 0 16000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_139
timestamp 0
transform 1 0 44000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_140
timestamp 0
transform 1 0 72000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_141
timestamp 0
transform 1 0 100000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_142
timestamp 0
transform 1 0 128000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_143
timestamp 0
transform 1 0 156000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_144
timestamp 0
transform 1 0 184000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_145
timestamp 0
transform 1 0 212000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_146
timestamp 0
transform 1 0 240000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_147
timestamp 0
transform 1 0 268000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_148
timestamp 0
transform 1 0 296000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_149
timestamp 0
transform 1 0 324000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_150
timestamp 0
transform 1 0 352000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_151
timestamp 0
transform 1 0 380000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_152
timestamp 0
transform 1 0 408000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_153
timestamp 0
transform 1 0 436000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_154
timestamp 0
transform 1 0 464000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_155
timestamp 0
transform 1 0 492000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_156
timestamp 0
transform 1 0 520000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_157
timestamp 0
transform 1 0 548000 0 1 205000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_158
timestamp 0
transform 1 0 16000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_159
timestamp 0
transform 1 0 44000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_160
timestamp 0
transform 1 0 72000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_161
timestamp 0
transform 1 0 100000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_162
timestamp 0
transform 1 0 128000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_163
timestamp 0
transform 1 0 156000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_164
timestamp 0
transform 1 0 184000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_165
timestamp 0
transform 1 0 212000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_166
timestamp 0
transform 1 0 240000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_167
timestamp 0
transform 1 0 268000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_168
timestamp 0
transform 1 0 296000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_169
timestamp 0
transform 1 0 324000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_170
timestamp 0
transform 1 0 352000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_171
timestamp 0
transform 1 0 380000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_172
timestamp 0
transform 1 0 408000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_173
timestamp 0
transform 1 0 436000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_174
timestamp 0
transform 1 0 464000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_175
timestamp 0
transform 1 0 492000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_176
timestamp 0
transform 1 0 520000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_177
timestamp 0
transform 1 0 548000 0 1 232000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_178
timestamp 0
transform 1 0 16000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_179
timestamp 0
transform 1 0 44000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_180
timestamp 0
transform 1 0 72000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_181
timestamp 0
transform 1 0 100000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_182
timestamp 0
transform 1 0 128000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_183
timestamp 0
transform 1 0 156000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_184
timestamp 0
transform 1 0 184000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_185
timestamp 0
transform 1 0 212000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_186
timestamp 0
transform 1 0 240000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_187
timestamp 0
transform 1 0 268000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_188
timestamp 0
transform 1 0 296000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_189
timestamp 0
transform 1 0 324000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_190
timestamp 0
transform 1 0 352000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_191
timestamp 0
transform 1 0 380000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_192
timestamp 0
transform 1 0 408000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_193
timestamp 0
transform 1 0 436000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_194
timestamp 0
transform 1 0 464000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_195
timestamp 0
transform 1 0 492000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_196
timestamp 0
transform 1 0 520000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_197
timestamp 0
transform 1 0 548000 0 1 259000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_198
timestamp 0
transform 1 0 16000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_199
timestamp 0
transform 1 0 44000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_200
timestamp 0
transform 1 0 72000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_201
timestamp 0
transform 1 0 100000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_202
timestamp 0
transform 1 0 128000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_203
timestamp 0
transform 1 0 156000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_204
timestamp 0
transform 1 0 184000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_205
timestamp 0
transform 1 0 212000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_206
timestamp 0
transform 1 0 240000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_207
timestamp 0
transform 1 0 268000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_208
timestamp 0
transform 1 0 296000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_209
timestamp 0
transform 1 0 324000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_210
timestamp 0
transform 1 0 352000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_211
timestamp 0
transform 1 0 380000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_212
timestamp 0
transform 1 0 408000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_213
timestamp 0
transform 1 0 436000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_214
timestamp 0
transform 1 0 464000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_215
timestamp 0
transform 1 0 492000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_216
timestamp 0
transform 1 0 520000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_217
timestamp 0
transform 1 0 548000 0 1 286000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_218
timestamp 0
transform 1 0 16000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_219
timestamp 0
transform 1 0 44000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_220
timestamp 0
transform 1 0 72000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_221
timestamp 0
transform 1 0 100000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_222
timestamp 0
transform 1 0 128000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_223
timestamp 0
transform 1 0 156000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_224
timestamp 0
transform 1 0 184000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_225
timestamp 0
transform 1 0 212000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_226
timestamp 0
transform 1 0 240000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_227
timestamp 0
transform 1 0 268000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_228
timestamp 0
transform 1 0 296000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_229
timestamp 0
transform 1 0 324000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_230
timestamp 0
transform 1 0 352000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_231
timestamp 0
transform 1 0 380000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_232
timestamp 0
transform 1 0 408000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_233
timestamp 0
transform 1 0 436000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_234
timestamp 0
transform 1 0 464000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_235
timestamp 0
transform 1 0 492000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_236
timestamp 0
transform 1 0 520000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_237
timestamp 0
transform 1 0 548000 0 1 313000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_238
timestamp 0
transform 1 0 16000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_239
timestamp 0
transform 1 0 44000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_240
timestamp 0
transform 1 0 72000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_241
timestamp 0
transform 1 0 100000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_242
timestamp 0
transform 1 0 128000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_243
timestamp 0
transform 1 0 156000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_244
timestamp 0
transform 1 0 184000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_245
timestamp 0
transform 1 0 212000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_246
timestamp 0
transform 1 0 240000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_247
timestamp 0
transform 1 0 268000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_248
timestamp 0
transform 1 0 296000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_249
timestamp 0
transform 1 0 324000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_250
timestamp 0
transform 1 0 352000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_251
timestamp 0
transform 1 0 380000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_252
timestamp 0
transform 1 0 408000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_253
timestamp 0
transform 1 0 436000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_254
timestamp 0
transform 1 0 464000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_255
timestamp 0
transform 1 0 492000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_256
timestamp 0
transform 1 0 520000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_257
timestamp 0
transform 1 0 548000 0 1 340000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_258
timestamp 0
transform 1 0 16000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_259
timestamp 0
transform 1 0 44000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_260
timestamp 0
transform 1 0 72000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_261
timestamp 0
transform 1 0 100000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_262
timestamp 0
transform 1 0 128000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_263
timestamp 0
transform 1 0 156000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_264
timestamp 0
transform 1 0 184000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_265
timestamp 0
transform 1 0 212000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_266
timestamp 0
transform 1 0 240000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_267
timestamp 0
transform 1 0 268000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_268
timestamp 0
transform 1 0 296000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_269
timestamp 0
transform 1 0 324000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_270
timestamp 0
transform 1 0 352000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_271
timestamp 0
transform 1 0 380000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_272
timestamp 0
transform 1 0 408000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_273
timestamp 0
transform 1 0 436000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_274
timestamp 0
transform 1 0 464000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_275
timestamp 0
transform 1 0 492000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_276
timestamp 0
transform 1 0 520000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_277
timestamp 0
transform 1 0 548000 0 1 367000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_278
timestamp 0
transform 1 0 16000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_279
timestamp 0
transform 1 0 44000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_280
timestamp 0
transform 1 0 72000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_281
timestamp 0
transform 1 0 100000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_282
timestamp 0
transform 1 0 128000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_283
timestamp 0
transform 1 0 156000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_284
timestamp 0
transform 1 0 184000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_285
timestamp 0
transform 1 0 212000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_286
timestamp 0
transform 1 0 240000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_287
timestamp 0
transform 1 0 268000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_288
timestamp 0
transform 1 0 296000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_289
timestamp 0
transform 1 0 324000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_290
timestamp 0
transform 1 0 352000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_291
timestamp 0
transform 1 0 380000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_292
timestamp 0
transform 1 0 408000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_293
timestamp 0
transform 1 0 436000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_294
timestamp 0
transform 1 0 464000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_295
timestamp 0
transform 1 0 492000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_296
timestamp 0
transform 1 0 520000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_297
timestamp 0
transform 1 0 548000 0 1 394000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_298
timestamp 0
transform 1 0 16000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_299
timestamp 0
transform 1 0 44000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_300
timestamp 0
transform 1 0 72000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_301
timestamp 0
transform 1 0 100000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_302
timestamp 0
transform 1 0 128000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_303
timestamp 0
transform 1 0 156000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_304
timestamp 0
transform 1 0 184000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_305
timestamp 0
transform 1 0 212000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_306
timestamp 0
transform 1 0 240000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_307
timestamp 0
transform 1 0 268000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_308
timestamp 0
transform 1 0 296000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_309
timestamp 0
transform 1 0 324000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_310
timestamp 0
transform 1 0 352000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_311
timestamp 0
transform 1 0 380000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_312
timestamp 0
transform 1 0 408000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_313
timestamp 0
transform 1 0 436000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_314
timestamp 0
transform 1 0 464000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_315
timestamp 0
transform 1 0 492000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_316
timestamp 0
transform 1 0 520000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_317
timestamp 0
transform 1 0 548000 0 1 421000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_318
timestamp 0
transform 1 0 16000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_319
timestamp 0
transform 1 0 44000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_320
timestamp 0
transform 1 0 72000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_321
timestamp 0
transform 1 0 100000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_322
timestamp 0
transform 1 0 128000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_323
timestamp 0
transform 1 0 156000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_324
timestamp 0
transform 1 0 184000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_325
timestamp 0
transform 1 0 212000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_326
timestamp 0
transform 1 0 240000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_327
timestamp 0
transform 1 0 268000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_328
timestamp 0
transform 1 0 296000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_329
timestamp 0
transform 1 0 324000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_330
timestamp 0
transform 1 0 352000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_331
timestamp 0
transform 1 0 380000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_332
timestamp 0
transform 1 0 408000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_333
timestamp 0
transform 1 0 436000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_334
timestamp 0
transform 1 0 464000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_335
timestamp 0
transform 1 0 492000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_336
timestamp 0
transform 1 0 520000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_337
timestamp 0
transform 1 0 548000 0 1 448000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_338
timestamp 0
transform 1 0 16000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_339
timestamp 0
transform 1 0 44000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_340
timestamp 0
transform 1 0 72000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_341
timestamp 0
transform 1 0 100000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_342
timestamp 0
transform 1 0 128000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_343
timestamp 0
transform 1 0 156000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_344
timestamp 0
transform 1 0 184000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_345
timestamp 0
transform 1 0 212000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_346
timestamp 0
transform 1 0 240000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_347
timestamp 0
transform 1 0 268000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_348
timestamp 0
transform 1 0 296000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_349
timestamp 0
transform 1 0 324000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_350
timestamp 0
transform 1 0 352000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_351
timestamp 0
transform 1 0 380000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_352
timestamp 0
transform 1 0 408000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_353
timestamp 0
transform 1 0 436000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_354
timestamp 0
transform 1 0 464000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_355
timestamp 0
transform 1 0 492000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_356
timestamp 0
transform 1 0 520000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_357
timestamp 0
transform 1 0 548000 0 1 475000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_358
timestamp 0
transform 1 0 16000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_359
timestamp 0
transform 1 0 44000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_360
timestamp 0
transform 1 0 72000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_361
timestamp 0
transform 1 0 100000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_362
timestamp 0
transform 1 0 128000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_363
timestamp 0
transform 1 0 156000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_364
timestamp 0
transform 1 0 184000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_365
timestamp 0
transform 1 0 212000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_366
timestamp 0
transform 1 0 240000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_367
timestamp 0
transform 1 0 268000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_368
timestamp 0
transform 1 0 296000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_369
timestamp 0
transform 1 0 324000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_370
timestamp 0
transform 1 0 352000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_371
timestamp 0
transform 1 0 380000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_372
timestamp 0
transform 1 0 408000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_373
timestamp 0
transform 1 0 436000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_374
timestamp 0
transform 1 0 464000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_375
timestamp 0
transform 1 0 492000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_376
timestamp 0
transform 1 0 520000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_377
timestamp 0
transform 1 0 548000 0 1 502000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_378
timestamp 0
transform 1 0 16000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_379
timestamp 0
transform 1 0 44000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_380
timestamp 0
transform 1 0 72000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_381
timestamp 0
transform 1 0 100000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_382
timestamp 0
transform 1 0 128000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_383
timestamp 0
transform 1 0 156000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_384
timestamp 0
transform 1 0 184000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_385
timestamp 0
transform 1 0 212000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_386
timestamp 0
transform 1 0 240000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_387
timestamp 0
transform 1 0 268000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_388
timestamp 0
transform 1 0 296000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_389
timestamp 0
transform 1 0 324000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_390
timestamp 0
transform 1 0 352000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_391
timestamp 0
transform 1 0 380000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_392
timestamp 0
transform 1 0 408000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_393
timestamp 0
transform 1 0 436000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_394
timestamp 0
transform 1 0 464000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_395
timestamp 0
transform 1 0 492000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_396
timestamp 0
transform 1 0 520000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_397
timestamp 0
transform 1 0 548000 0 1 529000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_398
timestamp 0
transform 1 0 16000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_399
timestamp 0
transform 1 0 44000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_400
timestamp 0
transform 1 0 72000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_401
timestamp 0
transform 1 0 100000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_402
timestamp 0
transform 1 0 128000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_403
timestamp 0
transform 1 0 156000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_404
timestamp 0
transform 1 0 184000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_405
timestamp 0
transform 1 0 212000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_406
timestamp 0
transform 1 0 240000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_407
timestamp 0
transform 1 0 268000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_408
timestamp 0
transform 1 0 296000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_409
timestamp 0
transform 1 0 324000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_410
timestamp 0
transform 1 0 352000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_411
timestamp 0
transform 1 0 380000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_412
timestamp 0
transform 1 0 408000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_413
timestamp 0
transform 1 0 436000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_414
timestamp 0
transform 1 0 464000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_415
timestamp 0
transform 1 0 492000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_416
timestamp 0
transform 1 0 520000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_417
timestamp 0
transform 1 0 548000 0 1 556000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_418
timestamp 0
transform 1 0 16000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_419
timestamp 0
transform 1 0 44000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_420
timestamp 0
transform 1 0 72000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_421
timestamp 0
transform 1 0 100000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_422
timestamp 0
transform 1 0 128000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_423
timestamp 0
transform 1 0 156000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_424
timestamp 0
transform 1 0 184000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_425
timestamp 0
transform 1 0 212000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_426
timestamp 0
transform 1 0 240000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_427
timestamp 0
transform 1 0 268000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_428
timestamp 0
transform 1 0 296000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_429
timestamp 0
transform 1 0 324000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_430
timestamp 0
transform 1 0 352000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_431
timestamp 0
transform 1 0 380000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_432
timestamp 0
transform 1 0 408000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_433
timestamp 0
transform 1 0 436000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_434
timestamp 0
transform 1 0 464000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_435
timestamp 0
transform 1 0 492000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_436
timestamp 0
transform 1 0 520000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_437
timestamp 0
transform 1 0 548000 0 1 583000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_438
timestamp 0
transform 1 0 16000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_439
timestamp 0
transform 1 0 44000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_440
timestamp 0
transform 1 0 72000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_441
timestamp 0
transform 1 0 100000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_442
timestamp 0
transform 1 0 128000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_443
timestamp 0
transform 1 0 156000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_444
timestamp 0
transform 1 0 184000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_445
timestamp 0
transform 1 0 212000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_446
timestamp 0
transform 1 0 240000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_447
timestamp 0
transform 1 0 268000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_448
timestamp 0
transform 1 0 296000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_449
timestamp 0
transform 1 0 324000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_450
timestamp 0
transform 1 0 352000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_451
timestamp 0
transform 1 0 380000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_452
timestamp 0
transform 1 0 408000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_453
timestamp 0
transform 1 0 436000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_454
timestamp 0
transform 1 0 464000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_455
timestamp 0
transform 1 0 492000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_456
timestamp 0
transform 1 0 520000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_457
timestamp 0
transform 1 0 548000 0 1 610000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_458
timestamp 0
transform 1 0 16000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_459
timestamp 0
transform 1 0 44000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_460
timestamp 0
transform 1 0 72000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_461
timestamp 0
transform 1 0 100000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_462
timestamp 0
transform 1 0 128000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_463
timestamp 0
transform 1 0 156000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_464
timestamp 0
transform 1 0 184000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_465
timestamp 0
transform 1 0 212000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_466
timestamp 0
transform 1 0 240000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_467
timestamp 0
transform 1 0 268000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_468
timestamp 0
transform 1 0 296000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_469
timestamp 0
transform 1 0 324000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_470
timestamp 0
transform 1 0 352000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_471
timestamp 0
transform 1 0 380000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_472
timestamp 0
transform 1 0 408000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_473
timestamp 0
transform 1 0 436000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_474
timestamp 0
transform 1 0 464000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_475
timestamp 0
transform 1 0 492000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_476
timestamp 0
transform 1 0 520000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_477
timestamp 0
transform 1 0 548000 0 1 637000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_478
timestamp 0
transform 1 0 16000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_479
timestamp 0
transform 1 0 44000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_480
timestamp 0
transform 1 0 72000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_481
timestamp 0
transform 1 0 100000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_482
timestamp 0
transform 1 0 128000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_483
timestamp 0
transform 1 0 156000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_484
timestamp 0
transform 1 0 184000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_485
timestamp 0
transform 1 0 212000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_486
timestamp 0
transform 1 0 240000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_487
timestamp 0
transform 1 0 268000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_488
timestamp 0
transform 1 0 296000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_489
timestamp 0
transform 1 0 324000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_490
timestamp 0
transform 1 0 352000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_491
timestamp 0
transform 1 0 380000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_492
timestamp 0
transform 1 0 408000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_493
timestamp 0
transform 1 0 436000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_494
timestamp 0
transform 1 0 464000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_495
timestamp 0
transform 1 0 492000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_496
timestamp 0
transform 1 0 520000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339501025136214612  scan_wrapper_339501025136214612_497
timestamp 0
transform 1 0 548000 0 1 664000
box 0 0 20000 20000
use scan_wrapper_339502597164499540  scan_wrapper_339502597164499540_4
timestamp 0
transform 1 0 184000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339732875283792466  scan_wrapper_339732875283792466_5
timestamp 0
transform 1 0 212000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339865743461974612  scan_wrapper_339865743461974612_6
timestamp 0
transform 1 0 240000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_339898704941023827  scan_wrapper_339898704941023827_7
timestamp 0
transform 1 0 268000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340218629792465491  scan_wrapper_340218629792465491_8
timestamp 0
transform 1 0 296000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340285391309374034  scan_wrapper_340285391309374034_10
timestamp 0
transform 1 0 352000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340318610245288530  scan_wrapper_340318610245288530_9
timestamp 0
transform 1 0 324000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340661930553246290  scan_wrapper_340661930553246290_11
timestamp 0
transform 1 0 380000 0 1 16000
box 0 0 20000 20000
use scan_wrapper_340805072482992722  scan_wrapper_340805072482992722_12
timestamp 0
transform 1 0 408000 0 1 16000
box 0 0 20000 20000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 41494 686000 42114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69494 686000 70114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 97494 686000 98114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 125494 686000 126114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 153494 686000 154114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181494 686000 182114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 209494 686000 210114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 237494 686000 238114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 265494 686000 266114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 293494 686000 294114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 321494 686000 322114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 349494 686000 350114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 377494 686000 378114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 405494 686000 406114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433494 686000 434114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 461494 686000 462114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 489494 686000 490114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 517494 686000 518114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545494 686000 546114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 573494 -7654 574114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 26241 592650 26861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 53241 592650 53861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 80241 592650 80861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107241 592650 107861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 134241 592650 134861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 161241 592650 161861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 188241 592650 188861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 215241 592650 215861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 242241 592650 242861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 269241 592650 269861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 296241 592650 296861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 323241 592650 323861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 350241 592650 350861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377241 592650 377861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 404241 592650 404861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 431241 592650 431861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 458241 592650 458861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 485241 592650 485861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512241 592650 512861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 539241 592650 539861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 566241 592650 566861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 593241 592650 593861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 620241 592650 620861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647241 592650 647861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 674241 592650 674861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 701241 592650 701861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 37994 686000 38614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 -7654 66614 41000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 686000 66614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 93994 686000 94614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 121994 686000 122614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149994 686000 150614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 177994 686000 178614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 205994 686000 206614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 233994 686000 234614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 261994 686000 262614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 289994 686000 290614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 317994 686000 318614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345994 686000 346614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 373994 686000 374614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401994 686000 402614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 429994 686000 430614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 457994 686000 458614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 485994 686000 486614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 513994 686000 514614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 541994 686000 542614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 569994 686000 570614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 22866 592650 23486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 49866 592650 50486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 76866 592650 77486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 130866 592650 131486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 157866 592650 158486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 184866 592650 185486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 211866 592650 212486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 238866 592650 239486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 265866 592650 266486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 292866 592650 293486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 319866 592650 320486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 346866 592650 347486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 400866 592650 401486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 427866 592650 428486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 454866 592650 455486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 481866 592650 482486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 508866 592650 509486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 535866 592650 536486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 562866 592650 563486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 589866 592650 590486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 616866 592650 617486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 670866 592650 671486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 697866 592650 698486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
