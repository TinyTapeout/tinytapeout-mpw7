VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_controller
  CLASS BLOCK ;
  FOREIGN scan_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 100.000 ;
  PIN active_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END active_select[0]
  PIN active_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 96.000 158.290 100.000 ;
    END
  END active_select[1]
  PIN active_select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 0.000 219.470 4.000 ;
    END
  END active_select[2]
  PIN active_select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 0.000 129.310 4.000 ;
    END
  END active_select[3]
  PIN active_select[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 96.000 42.370 100.000 ;
    END
  END active_select[4]
  PIN active_select[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END active_select[5]
  PIN active_select[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END active_select[6]
  PIN active_select[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 96.000 164.730 100.000 ;
    END
  END active_select[7]
  PIN active_select[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END active_select[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END clk
  PIN driver_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 96.000 0.510 100.000 ;
    END
  END driver_sel[0]
  PIN driver_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 96.000 122.870 100.000 ;
    END
  END driver_sel[1]
  PIN inputs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 0.000 164.730 4.000 ;
    END
  END inputs[0]
  PIN inputs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.810 0.000 203.370 4.000 ;
    END
  END inputs[1]
  PIN inputs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 96.000 213.030 100.000 ;
    END
  END inputs[2]
  PIN inputs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 96.000 229.130 100.000 ;
    END
  END inputs[3]
  PIN inputs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 30.340 230.000 31.540 ;
    END
  END inputs[4]
  PIN inputs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.540 4.000 24.740 ;
    END
  END inputs[5]
  PIN inputs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 96.000 58.470 100.000 ;
    END
  END inputs[6]
  PIN inputs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 40.540 230.000 41.740 ;
    END
  END inputs[7]
  PIN la_scan_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 0.000 145.410 4.000 ;
    END
  END la_scan_clk
  PIN la_scan_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 64.340 230.000 65.540 ;
    END
  END la_scan_data_in
  PIN la_scan_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 0.000 213.030 4.000 ;
    END
  END la_scan_data_out
  PIN la_scan_latch_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END la_scan_latch_en
  PIN la_scan_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 96.000 64.910 100.000 ;
    END
  END la_scan_select
  PIN oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 0.000 106.770 4.000 ;
    END
  END oeb[0]
  PIN oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 57.540 230.000 58.740 ;
    END
  END oeb[10]
  PIN oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 74.540 230.000 75.740 ;
    END
  END oeb[11]
  PIN oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 0.000 138.970 4.000 ;
    END
  END oeb[12]
  PIN oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 0.000 187.270 4.000 ;
    END
  END oeb[13]
  PIN oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 0.000 16.610 4.000 ;
    END
  END oeb[14]
  PIN oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 96.000 174.390 100.000 ;
    END
  END oeb[15]
  PIN oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 0.000 55.250 4.000 ;
    END
  END oeb[16]
  PIN oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 96.000 26.270 100.000 ;
    END
  END oeb[17]
  PIN oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 47.340 230.000 48.540 ;
    END
  END oeb[18]
  PIN oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END oeb[19]
  PIN oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 96.000 74.570 100.000 ;
    END
  END oeb[1]
  PIN oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 0.000 39.150 4.000 ;
    END
  END oeb[20]
  PIN oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END oeb[21]
  PIN oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930 96.000 190.490 100.000 ;
    END
  END oeb[22]
  PIN oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 96.000 32.710 100.000 ;
    END
  END oeb[23]
  PIN oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 0.000 97.110 4.000 ;
    END
  END oeb[24]
  PIN oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END oeb[25]
  PIN oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END oeb[26]
  PIN oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 96.000 132.530 100.000 ;
    END
  END oeb[27]
  PIN oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 0.000 196.930 4.000 ;
    END
  END oeb[28]
  PIN oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 0.000 229.130 4.000 ;
    END
  END oeb[29]
  PIN oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END oeb[2]
  PIN oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 96.000 16.610 100.000 ;
    END
  END oeb[30]
  PIN oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 96.000 116.430 100.000 ;
    END
  END oeb[31]
  PIN oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 96.000 148.630 100.000 ;
    END
  END oeb[32]
  PIN oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.740 4.000 17.940 ;
    END
  END oeb[33]
  PIN oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END oeb[34]
  PIN oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END oeb[35]
  PIN oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 96.000 138.970 100.000 ;
    END
  END oeb[36]
  PIN oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 96.000 180.830 100.000 ;
    END
  END oeb[37]
  PIN oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 96.000 222.690 100.000 ;
    END
  END oeb[3]
  PIN oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 96.000 100.330 100.000 ;
    END
  END oeb[4]
  PIN oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 96.000 10.170 100.000 ;
    END
  END oeb[5]
  PIN oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 0.000 6.950 4.000 ;
    END
  END oeb[6]
  PIN oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 91.540 230.000 92.740 ;
    END
  END oeb[7]
  PIN oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END oeb[8]
  PIN oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END oeb[9]
  PIN outputs[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 81.340 230.000 82.540 ;
    END
  END outputs[0]
  PIN outputs[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 0.000 171.170 4.000 ;
    END
  END outputs[1]
  PIN outputs[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 96.000 90.670 100.000 ;
    END
  END outputs[2]
  PIN outputs[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 13.340 230.000 14.540 ;
    END
  END outputs[3]
  PIN outputs[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 0.000 23.050 4.000 ;
    END
  END outputs[4]
  PIN outputs[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 0.000 48.810 4.000 ;
    END
  END outputs[5]
  PIN outputs[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 0.000 81.010 4.000 ;
    END
  END outputs[6]
  PIN outputs[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 23.540 230.000 24.740 ;
    END
  END outputs[7]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 0.000 90.670 4.000 ;
    END
  END ready
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 96.000 206.590 100.000 ;
    END
  END reset
  PIN scan_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 96.000 196.930 100.000 ;
    END
  END scan_clk
  PIN scan_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 96.000 84.230 100.000 ;
    END
  END scan_data_in
  PIN scan_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 96.000 106.770 100.000 ;
    END
  END scan_data_out
  PIN scan_latch_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 0.000 113.210 4.000 ;
    END
  END scan_latch_en
  PIN scan_select
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.740 4.000 51.940 ;
    END
  END scan_select
  PIN set_clk_div
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 96.000 48.810 100.000 ;
    END
  END set_clk_div
  PIN slow_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.000 3.140 230.000 4.340 ;
    END
  END slow_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.090 10.640 33.690 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.830 10.640 88.430 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.570 10.640 143.170 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.310 10.640 197.910 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 59.460 10.640 61.060 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.200 10.640 115.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.940 10.640 170.540 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.680 10.640 225.280 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 224.480 87.125 ;
      LAYER met1 ;
        RECT 0.070 9.220 229.010 87.280 ;
      LAYER met2 ;
        RECT 0.790 95.720 9.330 96.000 ;
        RECT 10.450 95.720 15.770 96.000 ;
        RECT 16.890 95.720 25.430 96.000 ;
        RECT 26.550 95.720 31.870 96.000 ;
        RECT 32.990 95.720 41.530 96.000 ;
        RECT 42.650 95.720 47.970 96.000 ;
        RECT 49.090 95.720 57.630 96.000 ;
        RECT 58.750 95.720 64.070 96.000 ;
        RECT 65.190 95.720 73.730 96.000 ;
        RECT 74.850 95.720 83.390 96.000 ;
        RECT 84.510 95.720 89.830 96.000 ;
        RECT 90.950 95.720 99.490 96.000 ;
        RECT 100.610 95.720 105.930 96.000 ;
        RECT 107.050 95.720 115.590 96.000 ;
        RECT 116.710 95.720 122.030 96.000 ;
        RECT 123.150 95.720 131.690 96.000 ;
        RECT 132.810 95.720 138.130 96.000 ;
        RECT 139.250 95.720 147.790 96.000 ;
        RECT 148.910 95.720 157.450 96.000 ;
        RECT 158.570 95.720 163.890 96.000 ;
        RECT 165.010 95.720 173.550 96.000 ;
        RECT 174.670 95.720 179.990 96.000 ;
        RECT 181.110 95.720 189.650 96.000 ;
        RECT 190.770 95.720 196.090 96.000 ;
        RECT 197.210 95.720 205.750 96.000 ;
        RECT 206.870 95.720 212.190 96.000 ;
        RECT 213.310 95.720 221.850 96.000 ;
        RECT 222.970 95.720 228.290 96.000 ;
        RECT 0.100 4.280 228.980 95.720 ;
        RECT 0.790 4.000 6.110 4.280 ;
        RECT 7.230 4.000 15.770 4.280 ;
        RECT 16.890 4.000 22.210 4.280 ;
        RECT 23.330 4.000 31.870 4.280 ;
        RECT 32.990 4.000 38.310 4.280 ;
        RECT 39.430 4.000 47.970 4.280 ;
        RECT 49.090 4.000 54.410 4.280 ;
        RECT 55.530 4.000 64.070 4.280 ;
        RECT 65.190 4.000 70.510 4.280 ;
        RECT 71.630 4.000 80.170 4.280 ;
        RECT 81.290 4.000 89.830 4.280 ;
        RECT 90.950 4.000 96.270 4.280 ;
        RECT 97.390 4.000 105.930 4.280 ;
        RECT 107.050 4.000 112.370 4.280 ;
        RECT 113.490 4.000 122.030 4.280 ;
        RECT 123.150 4.000 128.470 4.280 ;
        RECT 129.590 4.000 138.130 4.280 ;
        RECT 139.250 4.000 144.570 4.280 ;
        RECT 145.690 4.000 154.230 4.280 ;
        RECT 155.350 4.000 163.890 4.280 ;
        RECT 165.010 4.000 170.330 4.280 ;
        RECT 171.450 4.000 179.990 4.280 ;
        RECT 181.110 4.000 186.430 4.280 ;
        RECT 187.550 4.000 196.090 4.280 ;
        RECT 197.210 4.000 202.530 4.280 ;
        RECT 203.650 4.000 212.190 4.280 ;
        RECT 213.310 4.000 218.630 4.280 ;
        RECT 219.750 4.000 228.290 4.280 ;
      LAYER met3 ;
        RECT 4.400 94.540 226.010 95.705 ;
        RECT 4.000 93.140 226.010 94.540 ;
        RECT 4.000 91.140 225.600 93.140 ;
        RECT 4.000 86.340 226.010 91.140 ;
        RECT 4.400 84.340 226.010 86.340 ;
        RECT 4.000 82.940 226.010 84.340 ;
        RECT 4.000 80.940 225.600 82.940 ;
        RECT 4.000 76.140 226.010 80.940 ;
        RECT 4.400 74.140 225.600 76.140 ;
        RECT 4.000 69.340 226.010 74.140 ;
        RECT 4.400 67.340 226.010 69.340 ;
        RECT 4.000 65.940 226.010 67.340 ;
        RECT 4.000 63.940 225.600 65.940 ;
        RECT 4.000 59.140 226.010 63.940 ;
        RECT 4.400 57.140 225.600 59.140 ;
        RECT 4.000 52.340 226.010 57.140 ;
        RECT 4.400 50.340 226.010 52.340 ;
        RECT 4.000 48.940 226.010 50.340 ;
        RECT 4.000 46.940 225.600 48.940 ;
        RECT 4.000 42.140 226.010 46.940 ;
        RECT 4.400 40.140 225.600 42.140 ;
        RECT 4.000 35.340 226.010 40.140 ;
        RECT 4.400 33.340 226.010 35.340 ;
        RECT 4.000 31.940 226.010 33.340 ;
        RECT 4.000 29.940 225.600 31.940 ;
        RECT 4.000 25.140 226.010 29.940 ;
        RECT 4.400 23.140 225.600 25.140 ;
        RECT 4.000 18.340 226.010 23.140 ;
        RECT 4.400 16.340 226.010 18.340 ;
        RECT 4.000 14.940 226.010 16.340 ;
        RECT 4.000 12.940 225.600 14.940 ;
        RECT 4.000 8.140 226.010 12.940 ;
        RECT 4.400 6.140 226.010 8.140 ;
        RECT 4.000 4.740 226.010 6.140 ;
        RECT 4.000 3.590 225.600 4.740 ;
  END
END scan_controller
END LIBRARY

