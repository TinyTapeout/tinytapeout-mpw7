VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1
  CLASS BLOCK ;
  FOREIGN scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 96.000 96.970 100.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 96.000 0.370 100.000 ;
    END
  END latch_enable_out
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 87.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.640 96.990 87.280 ;
      LAYER met2 ;
        RECT 0.650 95.720 48.110 96.000 ;
        RECT 48.950 95.720 96.410 96.000 ;
        RECT 0.100 4.280 96.960 95.720 ;
        RECT 0.650 4.000 48.110 4.280 ;
        RECT 48.950 4.000 96.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 52.040 96.000 87.205 ;
        RECT 4.400 50.640 96.000 52.040 ;
        RECT 4.000 48.640 96.000 50.640 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 10.715 96.000 47.240 ;
      LAYER met4 ;
        RECT 17.775 10.640 19.150 87.280 ;
        RECT 21.550 10.640 33.970 87.280 ;
        RECT 36.370 10.640 48.800 87.280 ;
        RECT 51.200 10.640 63.625 87.280 ;
        RECT 66.025 10.640 78.455 87.280 ;
        RECT 80.855 10.640 88.945 87.280 ;
  END
END scan_wrapper_bc4d7220e4fdbf20a574d56ea112a8e1
END LIBRARY

